magic
tech scmos
magscale 1 2
timestamp 1656222261
<< metal1 >>
rect -66 1216 -2 1416
rect 2152 1404 2242 1416
rect 237 1337 252 1343
rect 436 1337 451 1343
rect 2109 1337 2156 1343
rect 621 1317 668 1323
rect 781 1317 796 1323
rect 1188 1317 1203 1323
rect 1357 1317 1372 1323
rect 2068 1317 2083 1323
rect 804 1277 819 1283
rect 1380 1277 1395 1283
rect 2045 1277 2060 1283
rect -66 1204 24 1216
rect -66 816 -2 1204
rect 61 1097 76 1103
rect 596 1097 611 1103
rect 1076 1097 1091 1103
rect 1261 1097 1308 1103
rect 1380 1097 1420 1103
rect 2013 1097 2083 1103
rect 2013 1084 2019 1097
rect 653 1077 668 1083
rect 836 1077 851 1083
rect 1133 1077 1148 1083
rect 1492 1077 1507 1083
rect 2178 1016 2242 1404
rect 2152 1004 2242 1016
rect 116 937 131 943
rect 420 937 435 943
rect 676 937 691 943
rect 852 937 867 943
rect 1357 937 1372 943
rect 1508 937 1523 943
rect 733 917 748 923
rect 909 917 972 923
rect 1549 917 1596 923
rect 1828 917 1843 923
rect -66 804 24 816
rect -66 416 -2 804
rect 84 697 131 703
rect 1140 697 1155 703
rect 1517 697 1548 703
rect 541 677 556 683
rect 1245 677 1260 683
rect 1517 677 1523 697
rect 1613 697 1635 703
rect 1613 684 1619 697
rect 2178 616 2242 1004
rect 2152 604 2242 616
rect 244 537 259 543
rect 964 537 979 543
rect 1181 537 1196 543
rect 669 517 716 523
rect 781 517 828 523
rect 1204 477 1219 483
rect -66 404 24 416
rect -66 16 -2 404
rect 765 297 780 303
rect 1092 297 1116 303
rect 1197 297 1228 303
rect 116 277 131 283
rect 468 277 483 283
rect 1197 277 1203 297
rect 1421 297 1436 303
rect 1485 297 1555 303
rect 1597 297 1612 303
rect 1549 284 1555 297
rect 1773 297 1788 303
rect 2004 297 2019 303
rect 1300 277 1315 283
rect 1380 277 1395 283
rect 1908 277 1923 283
rect 2178 216 2242 604
rect 2152 204 2242 216
rect 477 124 483 143
rect 1277 137 1292 143
rect 1364 137 1379 143
rect 1668 137 1683 143
rect 61 117 108 123
rect 484 117 499 123
rect 836 77 851 83
rect 2109 77 2124 83
rect -66 4 24 16
rect 2178 4 2242 204
<< m2contact >>
rect 316 1356 324 1364
rect 972 1356 980 1364
rect 1548 1356 1556 1364
rect 1884 1356 1892 1364
rect 12 1336 20 1344
rect 124 1336 132 1344
rect 140 1336 148 1344
rect 252 1336 260 1344
rect 332 1336 340 1344
rect 428 1336 436 1344
rect 508 1336 516 1344
rect 572 1336 580 1344
rect 636 1336 644 1344
rect 732 1336 740 1344
rect 748 1336 756 1344
rect 1004 1336 1012 1344
rect 1148 1336 1156 1344
rect 1244 1336 1252 1344
rect 1308 1336 1316 1344
rect 1324 1336 1332 1344
rect 1580 1336 1588 1344
rect 1852 1336 1860 1344
rect 2156 1336 2164 1344
rect 28 1316 36 1324
rect 60 1316 68 1324
rect 76 1316 84 1324
rect 108 1316 116 1324
rect 188 1316 196 1324
rect 268 1316 276 1324
rect 300 1316 308 1324
rect 364 1316 372 1324
rect 380 1316 388 1324
rect 412 1316 420 1324
rect 460 1316 468 1324
rect 492 1316 500 1324
rect 524 1316 532 1324
rect 556 1316 564 1324
rect 588 1316 596 1324
rect 668 1316 676 1324
rect 684 1316 692 1324
rect 796 1316 804 1324
rect 1068 1316 1076 1324
rect 1180 1316 1188 1324
rect 1260 1316 1268 1324
rect 1292 1316 1300 1324
rect 1372 1316 1380 1324
rect 1644 1316 1652 1324
rect 1788 1316 1796 1324
rect 2060 1316 2068 1324
rect 1100 1296 1108 1304
rect 1676 1296 1684 1304
rect 1756 1296 1764 1304
rect 796 1276 804 1284
rect 1372 1276 1380 1284
rect 2060 1276 2068 1284
rect 1100 1236 1108 1244
rect 1676 1236 1684 1244
rect 1756 1236 1764 1244
rect 76 1096 84 1104
rect 140 1096 148 1104
rect 172 1096 180 1104
rect 188 1096 196 1104
rect 220 1096 228 1104
rect 268 1096 276 1104
rect 300 1096 308 1104
rect 316 1096 324 1104
rect 348 1096 356 1104
rect 428 1096 436 1104
rect 508 1096 516 1104
rect 540 1096 548 1104
rect 588 1096 596 1104
rect 684 1096 692 1104
rect 716 1096 724 1104
rect 780 1096 788 1104
rect 860 1096 868 1104
rect 892 1096 900 1104
rect 956 1096 964 1104
rect 972 1096 980 1104
rect 1004 1096 1012 1104
rect 1068 1096 1076 1104
rect 1164 1096 1172 1104
rect 1196 1096 1204 1104
rect 1308 1096 1316 1104
rect 1324 1096 1332 1104
rect 1372 1096 1380 1104
rect 1420 1096 1428 1104
rect 1436 1096 1444 1104
rect 1516 1096 1524 1104
rect 1548 1096 1556 1104
rect 1580 1096 1588 1104
rect 1612 1096 1620 1104
rect 1644 1096 1652 1104
rect 1676 1096 1684 1104
rect 1740 1096 1748 1104
rect 1852 1096 1860 1104
rect 1964 1096 1972 1104
rect 12 1076 20 1084
rect 108 1076 116 1084
rect 124 1076 132 1084
rect 236 1076 244 1084
rect 252 1076 260 1084
rect 364 1076 372 1084
rect 380 1076 388 1084
rect 476 1076 484 1084
rect 492 1076 500 1084
rect 556 1076 564 1084
rect 668 1076 676 1084
rect 732 1076 740 1084
rect 828 1076 836 1084
rect 924 1076 932 1084
rect 1020 1076 1028 1084
rect 1036 1076 1044 1084
rect 1148 1076 1156 1084
rect 1228 1076 1236 1084
rect 1276 1076 1284 1084
rect 1372 1076 1380 1084
rect 1388 1076 1396 1084
rect 1484 1076 1492 1084
rect 1564 1076 1572 1084
rect 1628 1076 1636 1084
rect 1692 1076 1700 1084
rect 1788 1076 1796 1084
rect 1804 1076 1812 1084
rect 1900 1076 1908 1084
rect 1916 1076 1924 1084
rect 2012 1076 2020 1084
rect 2028 1076 2036 1084
rect 2124 1076 2132 1084
rect 908 1056 916 1064
rect 1212 1056 1220 1064
rect 188 956 196 964
rect 604 956 612 964
rect 1148 956 1156 964
rect 1372 956 1380 964
rect 1676 956 1684 964
rect 1948 956 1956 964
rect 12 936 20 944
rect 108 936 116 944
rect 204 936 212 944
rect 300 936 308 944
rect 316 936 324 944
rect 412 936 420 944
rect 492 936 500 944
rect 588 936 596 944
rect 668 936 676 944
rect 780 936 788 944
rect 844 936 852 944
rect 956 936 964 944
rect 1180 936 1188 944
rect 1372 936 1380 944
rect 1436 936 1444 944
rect 1500 936 1508 944
rect 1564 936 1572 944
rect 1660 936 1668 944
rect 1692 936 1700 944
rect 1772 936 1780 944
rect 1788 936 1796 944
rect 1884 936 1892 944
rect 1932 936 1940 944
rect 2012 936 2020 944
rect 2060 936 2068 944
rect 2124 936 2132 944
rect 60 916 68 924
rect 140 916 148 924
rect 172 916 180 924
rect 236 916 244 924
rect 252 916 260 924
rect 284 916 292 924
rect 364 916 372 924
rect 444 916 452 924
rect 476 916 484 924
rect 508 916 516 924
rect 540 916 548 924
rect 556 916 564 924
rect 620 916 628 924
rect 652 916 660 924
rect 748 916 756 924
rect 796 916 804 924
rect 828 916 836 924
rect 972 916 980 924
rect 1244 916 1252 924
rect 1324 916 1332 924
rect 1388 916 1396 924
rect 1420 916 1428 924
rect 1452 916 1460 924
rect 1484 916 1492 924
rect 1596 916 1604 924
rect 1612 916 1620 924
rect 1724 916 1732 924
rect 1740 916 1748 924
rect 1820 916 1828 924
rect 1900 916 1908 924
rect 1964 916 1972 924
rect 1996 916 2004 924
rect 2028 916 2036 924
rect 2076 916 2084 924
rect 2108 916 2116 924
rect 1276 896 1284 904
rect 988 876 996 884
rect 1276 836 1284 844
rect 1836 776 1844 784
rect 2124 736 2132 744
rect 1836 716 1844 724
rect 28 696 36 704
rect 60 696 68 704
rect 76 696 84 704
rect 188 696 196 704
rect 220 696 228 704
rect 252 696 260 704
rect 284 696 292 704
rect 332 696 340 704
rect 364 696 372 704
rect 396 696 404 704
rect 428 696 436 704
rect 492 696 500 704
rect 572 696 580 704
rect 604 696 612 704
rect 620 696 628 704
rect 652 696 660 704
rect 732 696 740 704
rect 796 696 804 704
rect 860 696 868 704
rect 892 696 900 704
rect 972 696 980 704
rect 1036 696 1044 704
rect 1068 696 1076 704
rect 1132 696 1140 704
rect 1212 696 1220 704
rect 1276 696 1284 704
rect 1308 696 1316 704
rect 1388 696 1396 704
rect 1452 696 1460 704
rect 1484 696 1492 704
rect 12 676 20 684
rect 76 676 84 684
rect 172 676 180 684
rect 236 676 244 684
rect 300 676 308 684
rect 316 676 324 684
rect 380 676 388 684
rect 444 676 452 684
rect 556 676 564 684
rect 668 676 676 684
rect 684 676 692 684
rect 780 676 788 684
rect 828 676 836 684
rect 908 676 916 684
rect 924 676 932 684
rect 1020 676 1028 684
rect 1084 676 1092 684
rect 1100 676 1108 684
rect 1196 676 1204 684
rect 1260 676 1268 684
rect 1324 676 1332 684
rect 1340 676 1348 684
rect 1436 676 1444 684
rect 1500 676 1508 684
rect 1548 696 1556 704
rect 1564 696 1572 704
rect 1740 696 1748 704
rect 1868 696 1876 704
rect 1612 676 1620 684
rect 1660 676 1668 684
rect 1692 676 1700 684
rect 1788 676 1796 684
rect 1932 676 1940 684
rect 844 656 852 664
rect 1260 656 1268 664
rect 1676 656 1684 664
rect 1964 656 1972 664
rect 316 556 324 564
rect 604 556 612 564
rect 956 556 964 564
rect 1372 556 1380 564
rect 1884 556 1892 564
rect 12 536 20 544
rect 124 536 132 544
rect 140 536 148 544
rect 236 536 244 544
rect 332 536 340 544
rect 428 536 436 544
rect 444 536 452 544
rect 540 536 548 544
rect 588 536 596 544
rect 620 536 628 544
rect 716 536 724 544
rect 732 536 740 544
rect 796 536 804 544
rect 892 536 900 544
rect 940 536 948 544
rect 956 536 964 544
rect 1068 536 1076 544
rect 1084 536 1092 544
rect 1196 536 1204 544
rect 1404 536 1412 544
rect 1548 536 1556 544
rect 1596 536 1604 544
rect 1692 536 1700 544
rect 1916 536 1924 544
rect 2060 536 2068 544
rect 2156 536 2164 544
rect 28 516 36 524
rect 60 516 68 524
rect 76 516 84 524
rect 108 516 116 524
rect 188 516 196 524
rect 268 516 276 524
rect 300 516 308 524
rect 364 516 372 524
rect 380 516 388 524
rect 412 516 420 524
rect 492 516 500 524
rect 556 516 564 524
rect 716 516 724 524
rect 748 516 756 524
rect 828 516 836 524
rect 844 516 852 524
rect 908 516 916 524
rect 1004 516 1012 524
rect 1020 516 1028 524
rect 1052 516 1060 524
rect 1132 516 1140 524
rect 1468 516 1476 524
rect 1580 516 1588 524
rect 1628 516 1636 524
rect 1644 516 1652 524
rect 1676 516 1684 524
rect 1980 516 1988 524
rect 2108 516 2116 524
rect 1500 496 1508 504
rect 2012 496 2020 504
rect 1196 476 1204 484
rect 1724 476 1732 484
rect 1500 436 1508 444
rect 2012 436 2020 444
rect 60 296 68 304
rect 140 296 148 304
rect 172 296 180 304
rect 188 296 196 304
rect 220 296 228 304
rect 300 296 308 304
rect 412 296 420 304
rect 492 296 500 304
rect 524 296 532 304
rect 540 296 548 304
rect 572 296 580 304
rect 652 296 660 304
rect 780 296 788 304
rect 844 296 852 304
rect 876 296 884 304
rect 908 296 916 304
rect 940 296 948 304
rect 1004 296 1012 304
rect 1068 296 1076 304
rect 1084 296 1092 304
rect 1116 296 1124 304
rect 1148 296 1156 304
rect 1180 296 1188 304
rect 12 276 20 284
rect 108 276 116 284
rect 236 276 244 284
rect 252 276 260 284
rect 348 276 356 284
rect 364 276 372 284
rect 460 276 468 284
rect 588 276 596 284
rect 604 276 612 284
rect 700 276 708 284
rect 716 276 724 284
rect 812 276 820 284
rect 828 276 836 284
rect 892 276 900 284
rect 972 276 980 284
rect 1020 276 1028 284
rect 1116 276 1124 284
rect 1132 276 1140 284
rect 1228 296 1236 304
rect 1244 296 1252 304
rect 1324 296 1332 304
rect 1356 296 1364 304
rect 1436 296 1444 304
rect 1612 296 1620 304
rect 1676 296 1684 304
rect 1708 296 1716 304
rect 1788 296 1796 304
rect 1852 296 1860 304
rect 1884 296 1892 304
rect 1948 296 1956 304
rect 1996 296 2004 304
rect 2076 296 2084 304
rect 2124 296 2132 304
rect 1292 276 1300 284
rect 1372 276 1380 284
rect 1436 276 1444 284
rect 1532 276 1540 284
rect 1548 276 1556 284
rect 1644 276 1652 284
rect 1660 276 1668 284
rect 1724 276 1732 284
rect 1820 276 1828 284
rect 1836 276 1844 284
rect 1900 276 1908 284
rect 1964 276 1972 284
rect 2060 276 2068 284
rect 2108 276 2116 284
rect 2156 276 2164 284
rect 956 256 964 264
rect 1372 256 1380 264
rect 1900 256 1908 264
rect 172 156 180 164
rect 252 156 260 164
rect 540 156 548 164
rect 1004 156 1012 164
rect 1356 156 1364 164
rect 1660 156 1668 164
rect 1948 156 1956 164
rect 12 136 20 144
rect 108 136 116 144
rect 156 136 164 144
rect 188 136 196 144
rect 268 136 276 144
rect 364 136 372 144
rect 380 136 388 144
rect 524 136 532 144
rect 556 136 564 144
rect 604 136 612 144
rect 700 136 708 144
rect 716 136 724 144
rect 764 136 772 144
rect 1036 136 1044 144
rect 1180 136 1188 144
rect 1292 136 1300 144
rect 1356 136 1364 144
rect 1420 136 1428 144
rect 1516 136 1524 144
rect 1532 136 1540 144
rect 1596 136 1604 144
rect 1660 136 1668 144
rect 1772 136 1780 144
rect 1916 136 1924 144
rect 108 116 116 124
rect 124 116 132 124
rect 204 116 212 124
rect 236 116 244 124
rect 300 116 308 124
rect 316 116 324 124
rect 348 116 356 124
rect 428 116 436 124
rect 476 116 484 124
rect 588 116 596 124
rect 652 116 660 124
rect 748 116 756 124
rect 780 116 788 124
rect 812 116 820 124
rect 1100 116 1108 124
rect 1228 116 1236 124
rect 1308 116 1316 124
rect 1340 116 1348 124
rect 1404 116 1412 124
rect 1468 116 1476 124
rect 1548 116 1556 124
rect 1580 116 1588 124
rect 1612 116 1620 124
rect 1644 116 1652 124
rect 1708 116 1716 124
rect 1724 116 1732 124
rect 1756 116 1764 124
rect 1852 116 1860 124
rect 1132 96 1140 104
rect 1820 96 1828 104
rect 828 76 836 84
rect 2124 76 2132 84
rect 1132 36 1140 44
rect 1820 36 1828 44
<< metal2 >>
rect 196 1397 220 1403
rect 260 1397 275 1403
rect 13 1344 19 1356
rect 13 1204 19 1336
rect 77 1324 83 1396
rect 109 1363 115 1396
rect 141 1363 147 1396
rect 109 1357 147 1363
rect 141 1344 147 1357
rect 29 1284 35 1316
rect 13 1084 19 1156
rect 45 1123 51 1156
rect 61 1124 67 1316
rect 45 1117 60 1123
rect 109 1104 115 1316
rect 125 1284 131 1336
rect 253 1324 259 1336
rect 269 1324 275 1397
rect 301 1377 339 1383
rect 301 1324 307 1377
rect 189 1244 195 1316
rect 125 1084 131 1116
rect 141 1104 147 1156
rect 109 1043 115 1076
rect 109 1037 124 1043
rect 13 964 19 1036
rect 13 944 19 956
rect 109 944 115 996
rect 125 923 131 956
rect 141 944 147 1076
rect 125 917 140 923
rect 29 704 35 876
rect 61 844 67 916
rect 61 723 67 796
rect 45 717 67 723
rect 45 684 51 717
rect 109 704 115 916
rect 157 884 163 1196
rect 189 1104 195 1156
rect 221 1104 227 1276
rect 269 1104 275 1196
rect 301 1104 307 1156
rect 317 1104 323 1356
rect 333 1344 339 1377
rect 429 1344 435 1356
rect 461 1324 467 1463
rect 493 1324 499 1356
rect 509 1344 515 1463
rect 525 1457 547 1463
rect 749 1457 771 1463
rect 365 1263 371 1316
rect 333 1257 371 1263
rect 173 964 179 1096
rect 189 1044 195 1096
rect 260 1077 275 1083
rect 189 923 195 956
rect 205 944 211 956
rect 237 943 243 1076
rect 269 1044 275 1077
rect 221 937 243 943
rect 180 917 195 923
rect 189 704 195 876
rect 221 803 227 937
rect 253 924 259 996
rect 301 944 307 1036
rect 333 1004 339 1257
rect 461 1244 467 1316
rect 509 1284 515 1336
rect 525 1324 531 1457
rect 573 1344 579 1356
rect 749 1344 755 1457
rect 973 1364 979 1463
rect 573 1324 579 1336
rect 637 1323 643 1336
rect 733 1324 739 1336
rect 596 1317 643 1323
rect 493 1277 508 1283
rect 349 1124 355 1236
rect 397 1204 403 1236
rect 429 1197 444 1203
rect 349 1104 355 1116
rect 365 1084 371 1156
rect 381 1084 387 1116
rect 429 1104 435 1197
rect 477 1084 483 1156
rect 493 1084 499 1277
rect 509 1104 515 1236
rect 372 997 419 1003
rect 413 944 419 997
rect 237 804 243 916
rect 212 797 227 803
rect 221 783 227 797
rect 221 777 243 783
rect 221 704 227 756
rect 61 683 67 696
rect 237 684 243 777
rect 61 677 76 683
rect 13 604 19 676
rect 13 544 19 596
rect 77 543 83 676
rect 109 604 115 636
rect 173 604 179 676
rect 141 544 147 596
rect 221 583 227 676
rect 253 603 259 696
rect 244 597 259 603
rect 180 577 227 583
rect 237 544 243 556
rect 77 537 99 543
rect 93 523 99 537
rect 93 517 108 523
rect 29 484 35 516
rect 61 404 67 516
rect 13 284 19 396
rect 61 304 67 356
rect 77 324 83 516
rect 125 484 131 536
rect 141 444 147 536
rect 189 404 195 516
rect 237 483 243 516
rect 253 484 259 597
rect 269 564 275 796
rect 285 704 291 716
rect 285 644 291 696
rect 301 684 307 936
rect 317 844 323 936
rect 477 924 483 956
rect 365 884 371 916
rect 340 877 355 883
rect 317 684 323 756
rect 333 704 339 716
rect 301 637 316 643
rect 301 623 307 637
rect 285 617 307 623
rect 285 524 291 617
rect 317 564 323 596
rect 333 564 339 676
rect 349 644 355 877
rect 413 803 419 916
rect 445 844 451 916
rect 404 797 419 803
rect 365 684 371 696
rect 381 684 387 756
rect 397 704 403 796
rect 493 764 499 936
rect 509 924 515 1096
rect 525 804 531 1316
rect 557 1303 563 1316
rect 589 1303 595 1316
rect 557 1297 595 1303
rect 541 1104 547 1116
rect 557 1084 563 1196
rect 669 1084 675 1316
rect 685 1284 691 1316
rect 797 1284 803 1316
rect 685 1104 691 1196
rect 717 1004 723 1096
rect 733 1084 739 1116
rect 781 1104 787 1156
rect 797 1124 803 1276
rect 1005 1244 1011 1336
rect 1069 1324 1075 1463
rect 1325 1457 1347 1463
rect 1101 1244 1107 1296
rect 1005 1124 1011 1156
rect 829 1084 835 1116
rect 861 1084 867 1096
rect 893 1084 899 1096
rect 909 1064 915 1116
rect 973 1104 979 1116
rect 1005 1104 1011 1116
rect 957 1084 963 1096
rect 1037 1084 1043 1116
rect 1069 1104 1075 1236
rect 1133 1204 1139 1356
rect 1149 1284 1155 1336
rect 1181 1223 1187 1316
rect 1197 1244 1203 1316
rect 1245 1284 1251 1336
rect 1261 1324 1267 1396
rect 1325 1344 1331 1457
rect 1277 1317 1292 1323
rect 1277 1303 1283 1317
rect 1261 1297 1283 1303
rect 1213 1263 1219 1276
rect 1261 1263 1267 1297
rect 1309 1284 1315 1336
rect 1213 1257 1267 1263
rect 1165 1217 1187 1223
rect 1165 1164 1171 1217
rect 1165 1104 1171 1156
rect 1021 1004 1027 1076
rect 1149 1004 1155 1076
rect 589 944 595 956
rect 605 923 611 956
rect 845 944 851 996
rect 1181 964 1187 1196
rect 1204 1097 1219 1103
rect 1213 1064 1219 1097
rect 1229 1084 1235 1196
rect 1245 964 1251 1236
rect 1341 1204 1347 1396
rect 1373 1284 1379 1316
rect 1581 1204 1587 1336
rect 1677 1244 1683 1296
rect 1757 1244 1763 1296
rect 1277 1084 1283 1156
rect 1325 1137 1379 1143
rect 1309 1104 1315 1116
rect 1325 1104 1331 1137
rect 1373 1104 1379 1137
rect 1389 1084 1395 1156
rect 1437 1104 1443 1196
rect 1748 1157 1772 1163
rect 1517 1104 1523 1156
rect 1581 1104 1587 1156
rect 1597 1137 1731 1143
rect 1549 1083 1555 1096
rect 1597 1084 1603 1137
rect 1725 1124 1731 1137
rect 1645 1104 1651 1116
rect 1549 1077 1564 1083
rect 1373 1004 1379 1076
rect 1613 1004 1619 1096
rect 1677 1063 1683 1096
rect 1693 1084 1699 1116
rect 1741 1104 1747 1156
rect 1805 1084 1811 1116
rect 1853 1104 1859 1336
rect 2157 1324 2163 1336
rect 2061 1284 2067 1316
rect 2061 1164 2067 1276
rect 1901 1084 1907 1156
rect 2125 1084 2131 1156
rect 1677 1057 1699 1063
rect 1380 957 1459 963
rect 628 937 668 943
rect 781 924 787 936
rect 957 924 963 936
rect 605 917 620 923
rect 429 604 435 696
rect 557 684 563 916
rect 653 884 659 916
rect 749 884 755 916
rect 797 903 803 916
rect 781 897 803 903
rect 781 804 787 897
rect 829 884 835 916
rect 973 884 979 916
rect 989 844 995 876
rect 589 697 604 703
rect 445 644 451 676
rect 573 644 579 696
rect 301 543 307 556
rect 301 537 323 543
rect 205 477 243 483
rect 109 284 115 316
rect 157 297 172 303
rect 141 284 147 296
rect 109 144 115 196
rect 157 144 163 297
rect 189 283 195 296
rect 173 277 195 283
rect 173 164 179 277
rect 205 204 211 477
rect 269 444 275 516
rect 301 484 307 516
rect 317 444 323 537
rect 349 543 355 596
rect 429 544 435 596
rect 541 544 547 596
rect 349 537 387 543
rect 333 484 339 536
rect 381 524 387 537
rect 365 463 371 516
rect 365 457 387 463
rect 381 444 387 457
rect 221 324 227 356
rect 221 304 227 316
rect 253 284 259 316
rect 301 304 307 356
rect 349 284 355 436
rect 413 404 419 516
rect 445 404 451 536
rect 493 484 499 516
rect 365 284 371 356
rect 413 304 419 356
rect 461 284 467 436
rect 557 404 563 516
rect 573 484 579 636
rect 589 544 595 697
rect 621 683 627 696
rect 653 684 659 696
rect 669 684 675 796
rect 733 704 739 756
rect 781 684 787 796
rect 605 677 627 683
rect 605 564 611 677
rect 797 644 803 696
rect 845 664 851 796
rect 893 724 899 756
rect 893 704 899 716
rect 861 684 867 696
rect 925 684 931 716
rect 973 704 979 756
rect 1021 684 1027 836
rect 1037 704 1043 796
rect 1069 704 1075 756
rect 1149 724 1155 956
rect 1181 764 1187 936
rect 1245 924 1251 956
rect 1277 844 1283 896
rect 1069 684 1075 696
rect 749 564 755 636
rect 717 544 723 556
rect 621 524 627 536
rect 733 524 739 536
rect 749 524 755 556
rect 893 544 899 596
rect 781 537 796 543
rect 717 444 723 516
rect 781 404 787 537
rect 829 484 835 516
rect 573 304 579 356
rect 589 324 595 396
rect 365 244 371 276
rect 493 244 499 296
rect 13 124 19 136
rect 189 124 195 136
rect 205 124 211 196
rect 356 157 387 163
rect 109 84 115 116
rect 221 84 227 156
rect 253 124 259 156
rect 237 103 243 116
rect 269 103 275 136
rect 349 124 355 156
rect 381 144 387 157
rect 365 124 371 136
rect 237 97 275 103
rect 301 84 307 116
rect 429 83 435 116
rect 493 103 499 156
rect 525 144 531 296
rect 541 164 547 296
rect 589 284 595 316
rect 605 284 611 356
rect 653 337 755 343
rect 653 304 659 337
rect 749 324 755 337
rect 701 284 707 316
rect 781 304 787 396
rect 813 284 819 316
rect 845 304 851 316
rect 477 97 499 103
rect 477 83 483 97
rect 429 77 483 83
rect 557 -17 563 136
rect 589 124 595 256
rect 877 244 883 296
rect 893 284 899 536
rect 909 524 915 676
rect 957 637 972 643
rect 957 564 963 637
rect 909 304 915 396
rect 941 323 947 536
rect 957 484 963 536
rect 1021 524 1027 636
rect 1085 604 1091 676
rect 1197 604 1203 676
rect 1069 544 1075 556
rect 1197 544 1203 556
rect 1213 543 1219 696
rect 1204 537 1219 543
rect 925 317 947 323
rect 605 144 611 156
rect 717 144 723 236
rect 605 124 611 136
rect 701 124 707 136
rect 733 123 739 196
rect 765 124 771 136
rect 781 124 787 156
rect 717 117 739 123
rect 653 44 659 116
rect 717 103 723 117
rect 756 117 764 123
rect 701 97 723 103
rect 701 44 707 97
rect 557 -23 579 -17
rect 733 -23 739 36
rect 781 23 787 76
rect 797 44 803 236
rect 813 84 819 116
rect 829 84 835 116
rect 909 44 915 116
rect 813 37 828 43
rect 813 23 819 37
rect 781 17 819 23
rect 925 -23 931 317
rect 948 297 963 303
rect 957 264 963 297
rect 989 283 995 476
rect 1005 403 1011 516
rect 1021 423 1027 476
rect 1053 444 1059 516
rect 1085 444 1091 536
rect 1245 484 1251 716
rect 1261 697 1276 703
rect 1261 684 1267 697
rect 1261 644 1267 656
rect 1220 477 1244 483
rect 1021 417 1043 423
rect 1005 397 1020 403
rect 1005 304 1011 356
rect 1021 284 1027 396
rect 1037 343 1043 417
rect 1037 337 1059 343
rect 1053 323 1059 337
rect 1053 317 1075 323
rect 1069 304 1075 317
rect 1085 304 1091 396
rect 1117 324 1123 436
rect 1124 297 1139 303
rect 1133 284 1139 297
rect 989 277 1011 283
rect 973 244 979 276
rect 1005 244 1011 277
rect 1117 263 1123 276
rect 1149 263 1155 296
rect 1117 257 1155 263
rect 1149 244 1155 257
rect 1005 44 1011 156
rect 1037 144 1043 236
rect 1044 37 1059 43
rect 1053 23 1059 37
rect 1053 17 1068 23
rect 1117 23 1123 156
rect 1149 124 1155 156
rect 1133 44 1139 96
rect 1165 44 1171 476
rect 1197 444 1203 476
rect 1293 423 1299 956
rect 1373 923 1379 936
rect 1373 917 1388 923
rect 1325 723 1331 916
rect 1421 884 1427 916
rect 1437 804 1443 936
rect 1453 924 1459 957
rect 1469 924 1475 956
rect 1501 944 1507 996
rect 1677 964 1683 996
rect 1693 944 1699 1057
rect 1485 844 1491 916
rect 1325 717 1340 723
rect 1453 723 1459 756
rect 1485 724 1491 756
rect 1517 724 1523 916
rect 1565 884 1571 936
rect 1597 823 1603 916
rect 1613 884 1619 916
rect 1613 844 1619 876
rect 1597 817 1635 823
rect 1453 717 1475 723
rect 1309 704 1315 716
rect 1341 684 1347 716
rect 1389 704 1395 716
rect 1453 644 1459 696
rect 1469 564 1475 717
rect 1485 704 1491 716
rect 1501 644 1507 676
rect 1373 484 1379 556
rect 1405 524 1411 536
rect 1469 484 1475 516
rect 1373 444 1379 476
rect 1501 444 1507 496
rect 1517 484 1523 716
rect 1549 704 1555 756
rect 1581 723 1587 756
rect 1565 717 1587 723
rect 1565 704 1571 717
rect 1613 644 1619 676
rect 1597 544 1603 596
rect 1293 417 1331 423
rect 1245 357 1260 363
rect 1229 324 1235 356
rect 1229 304 1235 316
rect 1245 304 1251 357
rect 1293 304 1299 356
rect 1188 297 1203 303
rect 1197 243 1203 297
rect 1197 237 1260 243
rect 1181 144 1187 196
rect 1293 163 1299 276
rect 1277 157 1299 163
rect 1181 124 1187 136
rect 1213 83 1219 116
rect 1229 103 1235 116
rect 1229 97 1251 103
rect 1245 83 1251 97
rect 1277 83 1283 157
rect 1309 143 1315 396
rect 1325 343 1331 417
rect 1549 404 1555 536
rect 1629 524 1635 817
rect 1661 804 1667 936
rect 1773 924 1779 936
rect 1693 917 1724 923
rect 1677 684 1683 756
rect 1693 684 1699 917
rect 1789 884 1795 936
rect 1885 924 1891 936
rect 1917 924 1923 1076
rect 2013 963 2019 1076
rect 2029 1044 2035 1076
rect 2029 1004 2035 1036
rect 1997 957 2019 963
rect 1741 704 1747 756
rect 1645 524 1651 636
rect 1588 517 1628 523
rect 1565 444 1571 516
rect 1629 484 1635 516
rect 1581 437 1596 443
rect 1581 423 1587 437
rect 1565 417 1587 423
rect 1325 337 1347 343
rect 1325 304 1331 316
rect 1341 183 1347 337
rect 1364 297 1379 303
rect 1373 284 1379 297
rect 1373 244 1379 256
rect 1325 177 1347 183
rect 1325 164 1331 177
rect 1341 157 1356 163
rect 1300 137 1315 143
rect 1293 124 1299 136
rect 1341 124 1347 157
rect 1213 77 1235 83
rect 1245 77 1283 83
rect 1229 43 1235 77
rect 1309 44 1315 116
rect 1357 84 1363 136
rect 1405 124 1411 356
rect 1421 283 1427 396
rect 1565 383 1571 417
rect 1549 377 1571 383
rect 1437 337 1475 343
rect 1437 304 1443 337
rect 1469 324 1475 337
rect 1549 324 1555 377
rect 1613 304 1619 396
rect 1645 284 1651 356
rect 1661 324 1667 676
rect 1677 644 1683 656
rect 1677 524 1683 596
rect 1693 544 1699 676
rect 1709 564 1715 636
rect 1684 457 1747 463
rect 1677 437 1724 443
rect 1677 404 1683 437
rect 1421 277 1436 283
rect 1421 144 1427 196
rect 1517 144 1523 236
rect 1533 163 1539 276
rect 1645 244 1651 276
rect 1677 244 1683 296
rect 1549 183 1555 196
rect 1549 177 1571 183
rect 1533 157 1555 163
rect 1421 84 1427 136
rect 1533 124 1539 136
rect 1549 124 1555 157
rect 1565 124 1571 177
rect 1597 164 1603 236
rect 1693 204 1699 316
rect 1709 304 1715 396
rect 1741 343 1747 457
rect 1725 337 1747 343
rect 1725 284 1731 337
rect 1773 304 1779 636
rect 1789 604 1795 676
rect 1805 463 1811 716
rect 1821 644 1827 916
rect 1901 844 1907 916
rect 1933 884 1939 936
rect 1949 923 1955 956
rect 1997 924 2003 957
rect 2013 924 2019 936
rect 2061 924 2067 936
rect 2109 924 2115 996
rect 2125 944 2131 1076
rect 1949 917 1964 923
rect 2020 917 2028 923
rect 2077 884 2083 916
rect 1837 724 1843 776
rect 1965 764 1971 836
rect 1869 704 1875 716
rect 1933 684 1939 756
rect 2125 744 2131 796
rect 1965 644 1971 656
rect 1821 604 1827 636
rect 1869 623 1875 636
rect 1869 617 1891 623
rect 1885 564 1891 617
rect 1981 564 1987 596
rect 1885 524 1891 556
rect 1789 457 1811 463
rect 1789 364 1795 457
rect 1805 343 1811 436
rect 1869 423 1875 436
rect 1837 417 1875 423
rect 1837 364 1843 417
rect 1805 337 1827 343
rect 1789 304 1795 316
rect 1821 303 1827 337
rect 1885 323 1891 516
rect 1917 484 1923 536
rect 1917 437 1932 443
rect 1869 317 1891 323
rect 1821 297 1852 303
rect 1821 284 1827 297
rect 1725 223 1731 276
rect 1725 217 1747 223
rect 1668 157 1683 163
rect 1597 144 1603 156
rect 1588 117 1603 123
rect 1373 77 1388 83
rect 1373 44 1379 77
rect 1469 83 1475 116
rect 1549 84 1555 116
rect 1469 77 1484 83
rect 1597 44 1603 117
rect 1661 123 1667 136
rect 1652 117 1667 123
rect 1677 44 1683 157
rect 1709 143 1715 156
rect 1693 137 1715 143
rect 1693 124 1699 137
rect 1725 124 1731 196
rect 1741 124 1747 217
rect 1757 164 1763 196
rect 1773 144 1779 236
rect 1805 164 1811 196
rect 1837 124 1843 276
rect 1853 124 1859 276
rect 1869 243 1875 317
rect 1885 263 1891 296
rect 1901 284 1907 396
rect 1917 284 1923 437
rect 1933 404 1939 436
rect 1981 404 1987 516
rect 1885 257 1900 263
rect 1933 263 1939 356
rect 1997 304 2003 476
rect 2013 444 2019 496
rect 2029 324 2035 596
rect 2045 524 2051 676
rect 2125 604 2131 736
rect 2061 544 2067 556
rect 2157 544 2163 756
rect 2157 364 2163 536
rect 2077 304 2083 316
rect 1949 284 1955 296
rect 1917 257 1939 263
rect 1869 237 1884 243
rect 1917 144 1923 257
rect 1949 164 1955 236
rect 1965 204 1971 276
rect 1709 44 1715 116
rect 1757 84 1763 116
rect 1821 44 1827 96
rect 1917 84 1923 116
rect 2029 44 2035 196
rect 2093 124 2099 356
rect 2109 284 2115 316
rect 2125 164 2131 296
rect 2125 84 2131 156
rect 1229 37 1244 43
rect 1325 37 1340 43
rect 1325 23 1331 37
rect 1117 17 1331 23
<< m3contact >>
rect 76 1396 84 1404
rect 108 1396 116 1404
rect 140 1396 148 1404
rect 188 1396 196 1404
rect 220 1396 228 1404
rect 252 1396 260 1404
rect 12 1356 20 1364
rect 28 1316 36 1324
rect 108 1316 116 1324
rect 28 1276 36 1284
rect 12 1196 20 1204
rect 12 1156 20 1164
rect 44 1156 52 1164
rect 60 1116 68 1124
rect 252 1316 260 1324
rect 124 1276 132 1284
rect 220 1276 228 1284
rect 188 1236 196 1244
rect 156 1196 164 1204
rect 140 1156 148 1164
rect 124 1116 132 1124
rect 76 1096 84 1104
rect 108 1096 116 1104
rect 140 1076 148 1084
rect 12 1036 20 1044
rect 124 1036 132 1044
rect 108 996 116 1004
rect 12 956 20 964
rect 124 956 132 964
rect 108 916 116 924
rect 140 936 148 944
rect 28 876 36 884
rect 60 836 68 844
rect 60 796 68 804
rect 188 1156 196 1164
rect 268 1196 276 1204
rect 300 1156 308 1164
rect 428 1356 436 1364
rect 492 1356 500 1364
rect 380 1316 388 1324
rect 412 1316 420 1324
rect 188 1036 196 1044
rect 172 956 180 964
rect 204 956 212 964
rect 268 1036 276 1044
rect 300 1036 308 1044
rect 252 996 260 1004
rect 156 876 164 884
rect 188 876 196 884
rect 204 796 212 804
rect 572 1356 580 1364
rect 972 1356 980 1364
rect 524 1316 532 1324
rect 572 1316 580 1324
rect 732 1316 740 1324
rect 348 1236 356 1244
rect 396 1236 404 1244
rect 460 1236 468 1244
rect 396 1196 404 1204
rect 364 1156 372 1164
rect 348 1116 356 1124
rect 380 1116 388 1124
rect 444 1196 452 1204
rect 476 1156 484 1164
rect 508 1276 516 1284
rect 508 1236 516 1244
rect 332 996 340 1004
rect 364 996 372 1004
rect 476 956 484 964
rect 284 916 292 924
rect 236 796 244 804
rect 268 796 276 804
rect 220 756 228 764
rect 76 696 84 704
rect 108 696 116 704
rect 12 676 20 684
rect 44 676 52 684
rect 220 676 228 684
rect 12 596 20 604
rect 108 636 116 644
rect 108 596 116 604
rect 140 596 148 604
rect 172 596 180 604
rect 172 576 180 584
rect 236 596 244 604
rect 236 556 244 564
rect 28 516 36 524
rect 28 476 36 484
rect 12 396 20 404
rect 60 396 68 404
rect 60 356 68 364
rect 124 476 132 484
rect 236 516 244 524
rect 140 436 148 444
rect 284 716 292 724
rect 412 916 420 924
rect 332 876 340 884
rect 316 836 324 844
rect 316 756 324 764
rect 332 716 340 724
rect 300 676 308 684
rect 332 676 340 684
rect 284 636 292 644
rect 316 636 324 644
rect 268 556 276 564
rect 316 596 324 604
rect 364 876 372 884
rect 396 796 404 804
rect 444 836 452 844
rect 380 756 388 764
rect 556 1196 564 1204
rect 540 1116 548 1124
rect 588 1096 596 1104
rect 684 1276 692 1284
rect 684 1196 692 1204
rect 780 1156 788 1164
rect 732 1116 740 1124
rect 1260 1396 1268 1404
rect 1132 1356 1140 1364
rect 1068 1316 1076 1324
rect 1004 1236 1012 1244
rect 1068 1236 1076 1244
rect 1004 1156 1012 1164
rect 796 1116 804 1124
rect 828 1116 836 1124
rect 908 1116 916 1124
rect 972 1116 980 1124
rect 1004 1116 1012 1124
rect 1036 1116 1044 1124
rect 732 1076 740 1084
rect 860 1076 868 1084
rect 892 1076 900 1084
rect 1196 1316 1204 1324
rect 1148 1276 1156 1284
rect 1340 1396 1348 1404
rect 1212 1276 1220 1284
rect 1244 1276 1252 1284
rect 1308 1276 1316 1284
rect 1196 1236 1204 1244
rect 1244 1236 1252 1244
rect 1132 1196 1140 1204
rect 1180 1196 1188 1204
rect 1228 1196 1236 1204
rect 1164 1156 1172 1164
rect 924 1076 932 1084
rect 956 1076 964 1084
rect 716 996 724 1004
rect 844 996 852 1004
rect 1020 996 1028 1004
rect 1148 996 1156 1004
rect 588 956 596 964
rect 540 916 548 924
rect 1548 1356 1556 1364
rect 1884 1356 1892 1364
rect 1372 1276 1380 1284
rect 1644 1316 1652 1324
rect 1788 1316 1796 1324
rect 1340 1196 1348 1204
rect 1436 1196 1444 1204
rect 1580 1196 1588 1204
rect 1276 1156 1284 1164
rect 1388 1156 1396 1164
rect 1308 1116 1316 1124
rect 1516 1156 1524 1164
rect 1580 1156 1588 1164
rect 1740 1156 1748 1164
rect 1772 1156 1780 1164
rect 1420 1096 1428 1104
rect 1388 1076 1396 1084
rect 1484 1076 1492 1084
rect 1644 1116 1652 1124
rect 1692 1116 1700 1124
rect 1724 1116 1732 1124
rect 1564 1076 1572 1084
rect 1596 1076 1604 1084
rect 1628 1076 1636 1084
rect 1804 1116 1812 1124
rect 2156 1316 2164 1324
rect 1900 1156 1908 1164
rect 2060 1156 2068 1164
rect 2124 1156 2132 1164
rect 1964 1096 1972 1104
rect 1788 1076 1796 1084
rect 1372 996 1380 1004
rect 1500 996 1508 1004
rect 1612 996 1620 1004
rect 1676 996 1684 1004
rect 1148 956 1156 964
rect 1180 956 1188 964
rect 1244 956 1252 964
rect 1292 956 1300 964
rect 620 936 628 944
rect 652 916 660 924
rect 780 916 788 924
rect 828 916 836 924
rect 956 916 964 924
rect 524 796 532 804
rect 492 756 500 764
rect 492 696 500 704
rect 364 676 372 684
rect 348 636 356 644
rect 652 876 660 884
rect 748 876 756 884
rect 828 876 836 884
rect 972 876 980 884
rect 988 836 996 844
rect 1020 836 1028 844
rect 668 796 676 804
rect 780 796 788 804
rect 844 796 852 804
rect 444 636 452 644
rect 572 636 580 644
rect 348 596 356 604
rect 428 596 436 604
rect 540 596 548 604
rect 300 556 308 564
rect 332 556 340 564
rect 284 516 292 524
rect 188 396 196 404
rect 76 316 84 324
rect 108 316 116 324
rect 12 276 20 284
rect 140 276 148 284
rect 108 196 116 204
rect 252 476 260 484
rect 300 476 308 484
rect 332 476 340 484
rect 268 436 276 444
rect 316 436 324 444
rect 348 436 356 444
rect 380 436 388 444
rect 220 356 228 364
rect 300 356 308 364
rect 220 316 228 324
rect 252 316 260 324
rect 492 476 500 484
rect 460 436 468 444
rect 412 396 420 404
rect 444 396 452 404
rect 364 356 372 364
rect 412 356 420 364
rect 732 756 740 764
rect 652 676 660 684
rect 684 676 692 684
rect 828 676 836 684
rect 892 756 900 764
rect 972 756 980 764
rect 892 716 900 724
rect 924 716 932 724
rect 1036 796 1044 804
rect 1068 756 1076 764
rect 1180 756 1188 764
rect 1148 716 1156 724
rect 1244 716 1252 724
rect 1132 696 1140 704
rect 860 676 868 684
rect 908 676 916 684
rect 1020 676 1028 684
rect 1068 676 1076 684
rect 1100 676 1108 684
rect 748 636 756 644
rect 796 636 804 644
rect 892 596 900 604
rect 716 556 724 564
rect 748 556 756 564
rect 620 516 628 524
rect 732 516 740 524
rect 572 476 580 484
rect 716 436 724 444
rect 844 516 852 524
rect 828 476 836 484
rect 556 396 564 404
rect 588 396 596 404
rect 780 396 788 404
rect 572 356 580 364
rect 604 356 612 364
rect 588 316 596 324
rect 236 276 244 284
rect 348 276 356 284
rect 364 236 372 244
rect 492 236 500 244
rect 204 196 212 204
rect 220 156 228 164
rect 348 156 356 164
rect 12 116 20 124
rect 124 116 132 124
rect 188 116 196 124
rect 252 116 260 124
rect 492 156 500 164
rect 316 116 324 124
rect 364 116 372 124
rect 476 116 484 124
rect 108 76 116 84
rect 220 76 228 84
rect 300 76 308 84
rect 700 316 708 324
rect 748 316 756 324
rect 812 316 820 324
rect 844 316 852 324
rect 716 276 724 284
rect 828 276 836 284
rect 588 256 596 264
rect 972 636 980 644
rect 1020 636 1028 644
rect 908 396 916 404
rect 1084 596 1092 604
rect 1196 596 1204 604
rect 1068 556 1076 564
rect 1196 556 1204 564
rect 956 476 964 484
rect 988 476 996 484
rect 716 236 724 244
rect 796 236 804 244
rect 876 236 884 244
rect 604 156 612 164
rect 732 196 740 204
rect 604 116 612 124
rect 700 116 708 124
rect 780 156 788 164
rect 764 116 772 124
rect 780 76 788 84
rect 652 36 660 44
rect 700 36 708 44
rect 732 36 740 44
rect 828 116 836 124
rect 908 116 916 124
rect 812 76 820 84
rect 796 36 804 44
rect 828 36 836 44
rect 908 36 916 44
rect 1020 476 1028 484
rect 1132 516 1140 524
rect 1260 636 1268 644
rect 1164 476 1172 484
rect 1212 476 1220 484
rect 1244 476 1252 484
rect 1052 436 1060 444
rect 1084 436 1092 444
rect 1116 436 1124 444
rect 1020 396 1028 404
rect 1004 356 1012 364
rect 1084 396 1092 404
rect 1116 316 1124 324
rect 972 236 980 244
rect 1004 236 1012 244
rect 1036 236 1044 244
rect 1148 236 1156 244
rect 1116 156 1124 164
rect 1148 156 1156 164
rect 1100 116 1108 124
rect 1004 36 1012 44
rect 1036 36 1044 44
rect 1068 16 1076 24
rect 1148 116 1156 124
rect 1196 436 1204 444
rect 1308 716 1316 724
rect 1420 876 1428 884
rect 1468 956 1476 964
rect 1468 916 1476 924
rect 1516 916 1524 924
rect 1484 836 1492 844
rect 1436 796 1444 804
rect 1452 756 1460 764
rect 1484 756 1492 764
rect 1340 716 1348 724
rect 1388 716 1396 724
rect 1596 916 1604 924
rect 1564 876 1572 884
rect 1612 876 1620 884
rect 1612 836 1620 844
rect 1548 756 1556 764
rect 1580 756 1588 764
rect 1324 676 1332 684
rect 1436 676 1444 684
rect 1452 636 1460 644
rect 1484 716 1492 724
rect 1516 716 1524 724
rect 1500 636 1508 644
rect 1468 556 1476 564
rect 1404 516 1412 524
rect 1372 476 1380 484
rect 1468 476 1476 484
rect 1612 636 1620 644
rect 1596 596 1604 604
rect 1516 476 1524 484
rect 1372 436 1380 444
rect 1308 396 1316 404
rect 1228 356 1236 364
rect 1228 316 1236 324
rect 1260 356 1268 364
rect 1292 356 1300 364
rect 1292 296 1300 304
rect 1260 236 1268 244
rect 1180 196 1188 204
rect 1180 116 1188 124
rect 1212 116 1220 124
rect 1660 796 1668 804
rect 1676 756 1684 764
rect 1740 916 1748 924
rect 1772 916 1780 924
rect 2028 1036 2036 1044
rect 2028 996 2036 1004
rect 2108 996 2116 1004
rect 1884 916 1892 924
rect 1916 916 1924 924
rect 1788 876 1796 884
rect 1740 756 1748 764
rect 1804 716 1812 724
rect 1676 676 1684 684
rect 1788 676 1796 684
rect 1644 636 1652 644
rect 1564 516 1572 524
rect 1628 476 1636 484
rect 1564 436 1572 444
rect 1596 436 1604 444
rect 1420 396 1428 404
rect 1548 396 1556 404
rect 1404 356 1412 364
rect 1324 316 1332 324
rect 1372 236 1380 244
rect 1324 156 1332 164
rect 1292 116 1300 124
rect 1164 36 1172 44
rect 1612 396 1620 404
rect 1468 316 1476 324
rect 1548 316 1556 324
rect 1644 356 1652 364
rect 1676 636 1684 644
rect 1676 596 1684 604
rect 1708 636 1716 644
rect 1772 636 1780 644
rect 1708 556 1716 564
rect 1724 476 1732 484
rect 1676 456 1684 464
rect 1724 436 1732 444
rect 1676 396 1684 404
rect 1708 396 1716 404
rect 1660 316 1668 324
rect 1692 316 1700 324
rect 1548 276 1556 284
rect 1660 276 1668 284
rect 1516 236 1524 244
rect 1420 196 1428 204
rect 1596 236 1604 244
rect 1644 236 1652 244
rect 1676 236 1684 244
rect 1548 196 1556 204
rect 1788 596 1796 604
rect 2012 916 2020 924
rect 2060 916 2068 924
rect 1932 876 1940 884
rect 2076 876 2084 884
rect 1900 836 1908 844
rect 1964 836 1972 844
rect 2124 796 2132 804
rect 1932 756 1940 764
rect 1964 756 1972 764
rect 1868 716 1876 724
rect 2156 756 2164 764
rect 2044 676 2052 684
rect 1820 636 1828 644
rect 1868 636 1876 644
rect 1964 636 1972 644
rect 1820 596 1828 604
rect 1980 596 1988 604
rect 2028 596 2036 604
rect 1980 556 1988 564
rect 1884 516 1892 524
rect 1804 436 1812 444
rect 1868 436 1876 444
rect 1788 356 1796 364
rect 1836 356 1844 364
rect 1788 316 1796 324
rect 1772 296 1780 304
rect 1916 476 1924 484
rect 1900 396 1908 404
rect 1852 276 1860 284
rect 1772 236 1780 244
rect 1692 196 1700 204
rect 1724 196 1732 204
rect 1596 156 1604 164
rect 1532 116 1540 124
rect 1564 116 1572 124
rect 1356 76 1364 84
rect 1388 76 1396 84
rect 1420 76 1428 84
rect 1484 76 1492 84
rect 1548 76 1556 84
rect 1612 116 1620 124
rect 1708 156 1716 164
rect 1756 196 1764 204
rect 1756 156 1764 164
rect 1804 196 1812 204
rect 1804 156 1812 164
rect 1932 436 1940 444
rect 1996 476 2004 484
rect 1932 396 1940 404
rect 1980 396 1988 404
rect 1932 356 1940 364
rect 1916 276 1924 284
rect 2124 596 2132 604
rect 2060 556 2068 564
rect 2044 516 2052 524
rect 2108 516 2116 524
rect 2092 356 2100 364
rect 2156 356 2164 364
rect 2028 316 2036 324
rect 2076 316 2084 324
rect 1948 276 1956 284
rect 2060 276 2068 284
rect 1884 236 1892 244
rect 1948 236 1956 244
rect 1964 196 1972 204
rect 2028 196 2036 204
rect 1692 116 1700 124
rect 1740 116 1748 124
rect 1836 116 1844 124
rect 1916 116 1924 124
rect 1756 76 1764 84
rect 1916 76 1924 84
rect 2108 316 2116 324
rect 2156 276 2164 284
rect 2124 156 2132 164
rect 2092 116 2100 124
rect 1244 36 1252 44
rect 1308 36 1316 44
rect 1340 36 1348 44
rect 1372 36 1380 44
rect 1596 36 1604 44
rect 1676 36 1684 44
rect 1708 36 1716 44
rect 2028 36 2036 44
<< metal3 >>
rect 74 1405 86 1406
rect 106 1405 118 1406
rect 74 1404 118 1405
rect 74 1396 76 1404
rect 84 1396 108 1404
rect 116 1396 118 1404
rect 74 1395 118 1396
rect 74 1394 86 1395
rect 106 1394 118 1395
rect 138 1405 150 1406
rect 186 1405 198 1406
rect 138 1404 198 1405
rect 138 1396 140 1404
rect 148 1396 188 1404
rect 196 1396 198 1404
rect 138 1395 198 1396
rect 138 1394 150 1395
rect 186 1394 198 1395
rect 218 1405 230 1406
rect 250 1405 262 1406
rect 218 1404 262 1405
rect 218 1396 220 1404
rect 228 1396 252 1404
rect 260 1396 262 1404
rect 218 1395 262 1396
rect 218 1394 230 1395
rect 250 1394 262 1395
rect 1258 1405 1270 1406
rect 1338 1405 1350 1406
rect 1258 1404 1350 1405
rect 1258 1396 1260 1404
rect 1268 1396 1340 1404
rect 1348 1396 1350 1404
rect 1258 1395 1350 1396
rect 1258 1394 1270 1395
rect 1338 1394 1350 1395
rect 10 1365 22 1366
rect 426 1365 438 1366
rect 10 1364 438 1365
rect 10 1356 12 1364
rect 20 1356 428 1364
rect 436 1356 438 1364
rect 10 1355 438 1356
rect 10 1354 22 1355
rect 426 1354 438 1355
rect 490 1365 502 1366
rect 570 1365 582 1366
rect 490 1364 582 1365
rect 490 1356 492 1364
rect 500 1356 572 1364
rect 580 1356 582 1364
rect 490 1355 582 1356
rect 490 1354 502 1355
rect 570 1354 582 1355
rect 970 1365 982 1366
rect 1130 1365 1142 1366
rect 1546 1365 1558 1366
rect 1882 1365 1894 1366
rect 970 1364 1894 1365
rect 970 1356 972 1364
rect 980 1356 1132 1364
rect 1140 1356 1548 1364
rect 1556 1356 1884 1364
rect 1892 1356 1894 1364
rect 970 1355 1894 1356
rect 970 1354 982 1355
rect 1130 1354 1142 1355
rect 1546 1354 1558 1355
rect 1882 1354 1894 1355
rect 26 1325 38 1326
rect 106 1325 118 1326
rect 26 1324 118 1325
rect 26 1316 28 1324
rect 36 1316 108 1324
rect 116 1316 118 1324
rect 26 1315 118 1316
rect 26 1314 38 1315
rect 106 1314 118 1315
rect 250 1325 262 1326
rect 378 1325 390 1326
rect 250 1324 390 1325
rect 250 1316 252 1324
rect 260 1316 380 1324
rect 388 1316 390 1324
rect 250 1315 390 1316
rect 250 1314 262 1315
rect 378 1314 390 1315
rect 410 1325 422 1326
rect 522 1325 534 1326
rect 410 1324 534 1325
rect 410 1316 412 1324
rect 420 1316 524 1324
rect 532 1316 534 1324
rect 410 1315 534 1316
rect 410 1314 422 1315
rect 522 1314 534 1315
rect 570 1325 582 1326
rect 730 1325 742 1326
rect 570 1324 742 1325
rect 570 1316 572 1324
rect 580 1316 732 1324
rect 740 1316 742 1324
rect 570 1315 742 1316
rect 570 1314 582 1315
rect 730 1314 742 1315
rect 1066 1325 1078 1326
rect 1194 1325 1206 1326
rect 1642 1325 1654 1326
rect 1786 1325 1798 1326
rect 1066 1324 1798 1325
rect 1066 1316 1068 1324
rect 1076 1316 1196 1324
rect 1204 1316 1644 1324
rect 1652 1316 1788 1324
rect 1796 1316 1798 1324
rect 1066 1315 1798 1316
rect 1066 1314 1078 1315
rect 1194 1314 1206 1315
rect 1642 1314 1654 1315
rect 1786 1314 1798 1315
rect 2154 1325 2166 1326
rect 2154 1324 2213 1325
rect 2154 1316 2156 1324
rect 2164 1316 2213 1324
rect 2154 1315 2213 1316
rect 2154 1314 2166 1315
rect -37 1285 -27 1305
rect 2203 1295 2213 1315
rect 26 1285 38 1286
rect -37 1284 38 1285
rect -37 1276 28 1284
rect 36 1276 38 1284
rect -37 1275 38 1276
rect 26 1274 38 1275
rect 122 1285 134 1286
rect 218 1285 230 1286
rect 506 1285 518 1286
rect 122 1284 518 1285
rect 122 1276 124 1284
rect 132 1276 220 1284
rect 228 1276 508 1284
rect 516 1276 518 1284
rect 122 1275 518 1276
rect 122 1274 134 1275
rect 218 1274 230 1275
rect 506 1274 518 1275
rect 682 1285 694 1286
rect 1146 1285 1158 1286
rect 1210 1285 1222 1286
rect 682 1284 1222 1285
rect 682 1276 684 1284
rect 692 1276 1148 1284
rect 1156 1276 1212 1284
rect 1220 1276 1222 1284
rect 682 1275 1222 1276
rect 682 1274 694 1275
rect 1146 1274 1158 1275
rect 1210 1274 1222 1275
rect 1242 1285 1254 1286
rect 1306 1285 1318 1286
rect 1370 1285 1382 1286
rect 1242 1284 1382 1285
rect 1242 1276 1244 1284
rect 1252 1276 1308 1284
rect 1316 1276 1372 1284
rect 1380 1276 1382 1284
rect 1242 1275 1382 1276
rect 1242 1274 1254 1275
rect 1306 1274 1318 1275
rect 1370 1274 1382 1275
rect 186 1245 198 1246
rect 346 1245 358 1246
rect 186 1244 358 1245
rect 186 1236 188 1244
rect 196 1236 348 1244
rect 356 1236 358 1244
rect 186 1235 358 1236
rect 186 1234 198 1235
rect 346 1234 358 1235
rect 394 1245 406 1246
rect 458 1245 470 1246
rect 506 1245 518 1246
rect 394 1244 518 1245
rect 394 1236 396 1244
rect 404 1236 460 1244
rect 468 1236 508 1244
rect 516 1236 518 1244
rect 394 1235 518 1236
rect 394 1234 406 1235
rect 458 1234 470 1235
rect 506 1234 518 1235
rect 1002 1245 1014 1246
rect 1066 1245 1078 1246
rect 1002 1244 1078 1245
rect 1002 1236 1004 1244
rect 1012 1236 1068 1244
rect 1076 1236 1078 1244
rect 1002 1235 1078 1236
rect 1002 1234 1014 1235
rect 1066 1234 1078 1235
rect 1194 1245 1206 1246
rect 1242 1245 1254 1246
rect 1194 1244 1254 1245
rect 1194 1236 1196 1244
rect 1204 1236 1244 1244
rect 1252 1236 1254 1244
rect 1194 1235 1254 1236
rect 1194 1234 1206 1235
rect 1242 1234 1254 1235
rect 10 1205 22 1206
rect 154 1205 166 1206
rect 10 1204 166 1205
rect 10 1196 12 1204
rect 20 1196 156 1204
rect 164 1196 166 1204
rect 10 1195 166 1196
rect 10 1194 22 1195
rect 154 1194 166 1195
rect 266 1205 278 1206
rect 394 1205 406 1206
rect 266 1204 406 1205
rect 266 1196 268 1204
rect 276 1196 396 1204
rect 404 1196 406 1204
rect 266 1195 406 1196
rect 266 1194 278 1195
rect 394 1194 406 1195
rect 442 1205 454 1206
rect 554 1205 566 1206
rect 682 1205 694 1206
rect 442 1204 694 1205
rect 442 1196 444 1204
rect 452 1196 556 1204
rect 564 1196 684 1204
rect 692 1196 694 1204
rect 442 1195 694 1196
rect 442 1194 454 1195
rect 554 1194 566 1195
rect 682 1194 694 1195
rect 1130 1205 1142 1206
rect 1178 1205 1190 1206
rect 1130 1204 1190 1205
rect 1130 1196 1132 1204
rect 1140 1196 1180 1204
rect 1188 1196 1190 1204
rect 1130 1195 1190 1196
rect 1130 1194 1142 1195
rect 1178 1194 1190 1195
rect 1226 1205 1238 1206
rect 1338 1205 1350 1206
rect 1226 1204 1350 1205
rect 1226 1196 1228 1204
rect 1236 1196 1340 1204
rect 1348 1196 1350 1204
rect 1226 1195 1350 1196
rect 1226 1194 1238 1195
rect 1338 1194 1350 1195
rect 1434 1205 1446 1206
rect 1578 1205 1590 1206
rect 1434 1204 1590 1205
rect 1434 1196 1436 1204
rect 1444 1196 1580 1204
rect 1588 1196 1590 1204
rect 1434 1195 1590 1196
rect 1434 1194 1446 1195
rect 1578 1194 1590 1195
rect 10 1165 22 1166
rect 42 1165 54 1166
rect 10 1164 54 1165
rect 10 1156 12 1164
rect 20 1156 44 1164
rect 52 1156 54 1164
rect 10 1155 54 1156
rect 10 1154 22 1155
rect 42 1154 54 1155
rect 138 1165 150 1166
rect 186 1165 198 1166
rect 138 1164 198 1165
rect 138 1156 140 1164
rect 148 1156 188 1164
rect 196 1156 198 1164
rect 138 1155 198 1156
rect 138 1154 150 1155
rect 186 1154 198 1155
rect 298 1165 310 1166
rect 362 1165 374 1166
rect 474 1165 486 1166
rect 298 1164 486 1165
rect 298 1156 300 1164
rect 308 1156 364 1164
rect 372 1156 476 1164
rect 484 1156 486 1164
rect 298 1155 486 1156
rect 298 1154 310 1155
rect 362 1154 374 1155
rect 474 1154 486 1155
rect 778 1165 790 1166
rect 1002 1165 1014 1166
rect 778 1164 1014 1165
rect 778 1156 780 1164
rect 788 1156 1004 1164
rect 1012 1156 1014 1164
rect 778 1155 1014 1156
rect 778 1154 790 1155
rect 1002 1154 1014 1155
rect 1162 1165 1174 1166
rect 1274 1165 1286 1166
rect 1162 1164 1286 1165
rect 1162 1156 1164 1164
rect 1172 1156 1276 1164
rect 1284 1156 1286 1164
rect 1162 1155 1286 1156
rect 1162 1154 1174 1155
rect 1274 1154 1286 1155
rect 1386 1165 1398 1166
rect 1514 1165 1526 1166
rect 1386 1164 1526 1165
rect 1386 1156 1388 1164
rect 1396 1156 1516 1164
rect 1524 1156 1526 1164
rect 1386 1155 1526 1156
rect 1386 1154 1398 1155
rect 1514 1154 1526 1155
rect 1578 1165 1590 1166
rect 1738 1165 1750 1166
rect 1578 1164 1750 1165
rect 1578 1156 1580 1164
rect 1588 1156 1740 1164
rect 1748 1156 1750 1164
rect 1578 1155 1750 1156
rect 1578 1154 1590 1155
rect 1738 1154 1750 1155
rect 1770 1165 1782 1166
rect 1898 1165 1910 1166
rect 1770 1164 1910 1165
rect 1770 1156 1772 1164
rect 1780 1156 1900 1164
rect 1908 1156 1910 1164
rect 1770 1155 1910 1156
rect 1770 1154 1782 1155
rect 1898 1154 1910 1155
rect 2058 1165 2070 1166
rect 2122 1165 2134 1166
rect 2058 1164 2134 1165
rect 2058 1156 2060 1164
rect 2068 1156 2124 1164
rect 2132 1156 2134 1164
rect 2058 1155 2134 1156
rect 2058 1154 2070 1155
rect 2122 1154 2134 1155
rect 58 1125 70 1126
rect 122 1125 134 1126
rect 58 1124 134 1125
rect 58 1116 60 1124
rect 68 1116 124 1124
rect 132 1116 134 1124
rect 58 1115 134 1116
rect 58 1114 70 1115
rect 122 1114 134 1115
rect 346 1125 358 1126
rect 378 1125 390 1126
rect 346 1124 390 1125
rect 346 1116 348 1124
rect 356 1116 380 1124
rect 388 1116 390 1124
rect 346 1115 390 1116
rect 346 1114 358 1115
rect 378 1114 390 1115
rect 538 1125 550 1126
rect 730 1125 742 1126
rect 538 1124 742 1125
rect 538 1116 540 1124
rect 548 1116 732 1124
rect 740 1116 742 1124
rect 538 1115 742 1116
rect 538 1114 550 1115
rect 730 1114 742 1115
rect 794 1125 806 1126
rect 826 1125 838 1126
rect 794 1124 838 1125
rect 794 1116 796 1124
rect 804 1116 828 1124
rect 836 1116 838 1124
rect 794 1115 838 1116
rect 794 1114 806 1115
rect 826 1114 838 1115
rect 906 1125 918 1126
rect 970 1125 982 1126
rect 906 1124 982 1125
rect 906 1116 908 1124
rect 916 1116 972 1124
rect 980 1116 982 1124
rect 906 1115 982 1116
rect 906 1114 918 1115
rect 970 1114 982 1115
rect 1002 1125 1014 1126
rect 1034 1125 1046 1126
rect 1002 1124 1046 1125
rect 1002 1116 1004 1124
rect 1012 1116 1036 1124
rect 1044 1116 1046 1124
rect 1002 1115 1046 1116
rect 1002 1114 1014 1115
rect 1034 1114 1046 1115
rect 1306 1125 1318 1126
rect 1642 1125 1654 1126
rect 1690 1125 1702 1126
rect 1306 1124 1702 1125
rect 1306 1116 1308 1124
rect 1316 1116 1644 1124
rect 1652 1116 1692 1124
rect 1700 1116 1702 1124
rect 1306 1115 1702 1116
rect 1306 1114 1318 1115
rect 1642 1114 1654 1115
rect 1690 1114 1702 1115
rect 1722 1125 1734 1126
rect 1802 1125 1814 1126
rect 1722 1124 1814 1125
rect 1722 1116 1724 1124
rect 1732 1116 1804 1124
rect 1812 1116 1814 1124
rect 1722 1115 1814 1116
rect 1722 1114 1734 1115
rect 1802 1114 1814 1115
rect 74 1104 86 1106
rect 74 1096 76 1104
rect 84 1096 86 1104
rect 74 1094 86 1096
rect 106 1104 118 1106
rect 106 1096 108 1104
rect 116 1096 118 1104
rect 106 1094 118 1096
rect 586 1104 598 1106
rect 586 1096 588 1104
rect 596 1096 598 1104
rect 586 1094 598 1096
rect 1418 1104 1430 1106
rect 1418 1096 1420 1104
rect 1428 1096 1430 1104
rect 1418 1094 1430 1096
rect 1962 1104 1974 1106
rect 1962 1096 1964 1104
rect 1972 1096 1974 1104
rect 1962 1094 1974 1096
rect 10 1045 22 1046
rect 75 1045 85 1094
rect 107 1085 117 1094
rect 138 1085 150 1086
rect 107 1084 150 1085
rect 107 1076 140 1084
rect 148 1076 150 1084
rect 107 1075 150 1076
rect 587 1085 597 1094
rect 730 1085 742 1086
rect 858 1085 870 1086
rect 587 1075 629 1085
rect 138 1074 150 1075
rect 10 1044 85 1045
rect 10 1036 12 1044
rect 20 1036 85 1044
rect 10 1035 85 1036
rect 122 1045 134 1046
rect 186 1045 198 1046
rect 122 1044 198 1045
rect 122 1036 124 1044
rect 132 1036 188 1044
rect 196 1036 198 1044
rect 122 1035 198 1036
rect 10 1034 22 1035
rect 122 1034 134 1035
rect 186 1034 198 1035
rect 266 1045 278 1046
rect 298 1045 310 1046
rect 266 1044 310 1045
rect 266 1036 268 1044
rect 276 1036 300 1044
rect 308 1036 310 1044
rect 266 1035 310 1036
rect 619 1045 629 1075
rect 730 1084 870 1085
rect 730 1076 732 1084
rect 740 1076 860 1084
rect 868 1076 870 1084
rect 730 1075 870 1076
rect 730 1074 742 1075
rect 858 1074 870 1075
rect 890 1085 902 1086
rect 922 1085 934 1086
rect 890 1084 934 1085
rect 890 1076 892 1084
rect 900 1076 924 1084
rect 932 1076 934 1084
rect 890 1075 934 1076
rect 890 1074 902 1075
rect 922 1074 934 1075
rect 954 1085 966 1086
rect 1386 1085 1398 1086
rect 954 1084 1398 1085
rect 954 1076 956 1084
rect 964 1076 1388 1084
rect 1396 1076 1398 1084
rect 954 1075 1398 1076
rect 1419 1085 1429 1094
rect 1482 1085 1494 1086
rect 1419 1084 1494 1085
rect 1419 1076 1484 1084
rect 1492 1076 1494 1084
rect 1419 1075 1494 1076
rect 954 1074 966 1075
rect 1386 1074 1398 1075
rect 1482 1074 1494 1075
rect 1562 1085 1574 1086
rect 1594 1085 1606 1086
rect 1562 1084 1606 1085
rect 1562 1076 1564 1084
rect 1572 1076 1596 1084
rect 1604 1076 1606 1084
rect 1562 1075 1606 1076
rect 1562 1074 1574 1075
rect 1594 1074 1606 1075
rect 1626 1085 1638 1086
rect 1786 1085 1798 1086
rect 1963 1085 1973 1094
rect 1626 1084 1973 1085
rect 1626 1076 1628 1084
rect 1636 1076 1788 1084
rect 1796 1076 1973 1084
rect 1626 1075 1973 1076
rect 1626 1074 1638 1075
rect 1786 1074 1798 1075
rect 2026 1045 2038 1046
rect 619 1044 2038 1045
rect 619 1036 2028 1044
rect 2036 1036 2038 1044
rect 619 1035 2038 1036
rect 266 1034 278 1035
rect 298 1034 310 1035
rect 2026 1034 2038 1035
rect 106 1005 118 1006
rect 250 1005 262 1006
rect 106 1004 262 1005
rect 106 996 108 1004
rect 116 996 252 1004
rect 260 996 262 1004
rect 106 995 262 996
rect 106 994 118 995
rect 250 994 262 995
rect 330 1005 342 1006
rect 362 1005 374 1006
rect 330 1004 374 1005
rect 330 996 332 1004
rect 340 996 364 1004
rect 372 996 374 1004
rect 330 995 374 996
rect 330 994 342 995
rect 362 994 374 995
rect 714 1005 726 1006
rect 842 1005 854 1006
rect 714 1004 854 1005
rect 714 996 716 1004
rect 724 996 844 1004
rect 852 996 854 1004
rect 714 995 854 996
rect 714 994 726 995
rect 842 994 854 995
rect 1018 1005 1030 1006
rect 1146 1005 1158 1006
rect 1370 1005 1382 1006
rect 1498 1005 1510 1006
rect 1018 1004 1510 1005
rect 1018 996 1020 1004
rect 1028 996 1148 1004
rect 1156 996 1372 1004
rect 1380 996 1500 1004
rect 1508 996 1510 1004
rect 1018 995 1510 996
rect 1018 994 1030 995
rect 1146 994 1158 995
rect 1370 994 1382 995
rect 1498 994 1510 995
rect 1610 1005 1622 1006
rect 1674 1005 1686 1006
rect 1610 1004 1686 1005
rect 1610 996 1612 1004
rect 1620 996 1676 1004
rect 1684 996 1686 1004
rect 1610 995 1686 996
rect 1610 994 1622 995
rect 1674 994 1686 995
rect 2026 1005 2038 1006
rect 2106 1005 2118 1006
rect 2026 1004 2118 1005
rect 2026 996 2028 1004
rect 2036 996 2108 1004
rect 2116 996 2118 1004
rect 2026 995 2118 996
rect 2026 994 2038 995
rect 2106 994 2118 995
rect 10 965 22 966
rect 122 965 134 966
rect 10 964 134 965
rect 10 956 12 964
rect 20 956 124 964
rect 132 956 134 964
rect 10 955 134 956
rect 10 954 22 955
rect 122 954 134 955
rect 170 965 182 966
rect 202 965 214 966
rect 170 964 214 965
rect 170 956 172 964
rect 180 956 204 964
rect 212 956 214 964
rect 170 955 214 956
rect 170 954 182 955
rect 202 954 214 955
rect 474 965 486 966
rect 586 965 598 966
rect 474 964 598 965
rect 474 956 476 964
rect 484 956 588 964
rect 596 956 598 964
rect 474 955 598 956
rect 474 954 486 955
rect 586 954 598 955
rect 1146 965 1158 966
rect 1178 965 1190 966
rect 1146 964 1190 965
rect 1146 956 1148 964
rect 1156 956 1180 964
rect 1188 956 1190 964
rect 1146 955 1190 956
rect 1146 954 1158 955
rect 1178 954 1190 955
rect 1242 965 1254 966
rect 1290 965 1302 966
rect 1466 965 1478 966
rect 1242 964 1478 965
rect 1242 956 1244 964
rect 1252 956 1292 964
rect 1300 956 1468 964
rect 1476 956 1478 964
rect 1242 955 1478 956
rect 1242 954 1254 955
rect 1290 954 1302 955
rect 1466 954 1478 955
rect 138 944 150 946
rect 138 936 140 944
rect 148 936 150 944
rect 138 934 150 936
rect 618 944 630 946
rect 618 936 620 944
rect 628 936 630 944
rect 618 934 630 936
rect 106 925 118 926
rect 139 925 149 934
rect -37 885 -27 925
rect 106 924 149 925
rect 106 916 108 924
rect 116 916 149 924
rect 106 915 149 916
rect 282 925 294 926
rect 410 925 422 926
rect 282 924 422 925
rect 282 916 284 924
rect 292 916 412 924
rect 420 916 422 924
rect 282 915 422 916
rect 106 914 118 915
rect 282 914 294 915
rect 410 914 422 915
rect 538 925 550 926
rect 619 925 629 934
rect 538 924 629 925
rect 538 916 540 924
rect 548 916 629 924
rect 538 915 629 916
rect 650 925 662 926
rect 778 925 790 926
rect 650 924 790 925
rect 650 916 652 924
rect 660 916 780 924
rect 788 916 790 924
rect 650 915 790 916
rect 538 914 550 915
rect 650 914 662 915
rect 778 914 790 915
rect 826 925 838 926
rect 954 925 966 926
rect 826 924 966 925
rect 826 916 828 924
rect 836 916 956 924
rect 964 916 966 924
rect 826 915 966 916
rect 826 914 838 915
rect 954 914 966 915
rect 1466 925 1478 926
rect 1514 925 1526 926
rect 1466 924 1526 925
rect 1466 916 1468 924
rect 1476 916 1516 924
rect 1524 916 1526 924
rect 1466 915 1526 916
rect 1466 914 1478 915
rect 1514 914 1526 915
rect 1594 925 1606 926
rect 1738 925 1750 926
rect 1594 924 1750 925
rect 1594 916 1596 924
rect 1604 916 1740 924
rect 1748 916 1750 924
rect 1594 915 1750 916
rect 1594 914 1606 915
rect 1738 914 1750 915
rect 1770 925 1782 926
rect 1882 925 1894 926
rect 1914 925 1926 926
rect 2010 925 2022 926
rect 1770 924 2022 925
rect 1770 916 1772 924
rect 1780 916 1884 924
rect 1892 916 1916 924
rect 1924 916 2012 924
rect 2020 916 2022 924
rect 1770 915 2022 916
rect 1770 914 1782 915
rect 1882 914 1894 915
rect 1914 914 1926 915
rect 2010 914 2022 915
rect 2058 925 2070 926
rect 2058 924 2213 925
rect 2058 916 2060 924
rect 2068 916 2213 924
rect 2058 915 2213 916
rect 2058 914 2070 915
rect 2203 895 2213 915
rect 26 885 38 886
rect 154 885 166 886
rect -37 884 166 885
rect -37 876 28 884
rect 36 876 156 884
rect 164 876 166 884
rect -37 875 166 876
rect 26 874 38 875
rect 154 874 166 875
rect 186 885 198 886
rect 330 885 342 886
rect 186 884 342 885
rect 186 876 188 884
rect 196 876 332 884
rect 340 876 342 884
rect 186 875 342 876
rect 186 874 198 875
rect 330 874 342 875
rect 362 885 374 886
rect 650 885 662 886
rect 362 884 662 885
rect 362 876 364 884
rect 372 876 652 884
rect 660 876 662 884
rect 362 875 662 876
rect 362 874 374 875
rect 650 874 662 875
rect 746 885 758 886
rect 826 885 838 886
rect 746 884 838 885
rect 746 876 748 884
rect 756 876 828 884
rect 836 876 838 884
rect 746 875 838 876
rect 746 874 758 875
rect 826 874 838 875
rect 970 885 982 886
rect 1418 885 1430 886
rect 1562 885 1574 886
rect 970 884 1574 885
rect 970 876 972 884
rect 980 876 1420 884
rect 1428 876 1564 884
rect 1572 876 1574 884
rect 970 875 1574 876
rect 970 874 982 875
rect 1418 874 1430 875
rect 1562 874 1574 875
rect 1610 885 1622 886
rect 1786 885 1798 886
rect 1610 884 1798 885
rect 1610 876 1612 884
rect 1620 876 1788 884
rect 1796 876 1798 884
rect 1610 875 1798 876
rect 1610 874 1622 875
rect 1786 874 1798 875
rect 1930 885 1942 886
rect 2074 885 2086 886
rect 1930 884 2086 885
rect 1930 876 1932 884
rect 1940 876 2076 884
rect 2084 876 2086 884
rect 1930 875 2086 876
rect 1930 874 1942 875
rect 2074 874 2086 875
rect 58 845 70 846
rect 314 845 326 846
rect 442 845 454 846
rect 58 844 454 845
rect 58 836 60 844
rect 68 836 316 844
rect 324 836 444 844
rect 452 836 454 844
rect 58 835 454 836
rect 58 834 70 835
rect 314 834 326 835
rect 442 834 454 835
rect 986 845 998 846
rect 1018 845 1030 846
rect 986 844 1030 845
rect 986 836 988 844
rect 996 836 1020 844
rect 1028 836 1030 844
rect 986 835 1030 836
rect 986 834 998 835
rect 1018 834 1030 835
rect 1482 845 1494 846
rect 1610 845 1622 846
rect 1482 844 1622 845
rect 1482 836 1484 844
rect 1492 836 1612 844
rect 1620 836 1622 844
rect 1482 835 1622 836
rect 1482 834 1494 835
rect 1610 834 1622 835
rect 1898 845 1910 846
rect 1962 845 1974 846
rect 1898 844 1974 845
rect 1898 836 1900 844
rect 1908 836 1964 844
rect 1972 836 1974 844
rect 1898 835 1974 836
rect 1898 834 1910 835
rect 1962 834 1974 835
rect 58 805 70 806
rect 202 805 214 806
rect 58 804 214 805
rect 58 796 60 804
rect 68 796 204 804
rect 212 796 214 804
rect 58 795 214 796
rect 58 794 70 795
rect 202 794 214 795
rect 234 805 246 806
rect 266 805 278 806
rect 234 804 278 805
rect 234 796 236 804
rect 244 796 268 804
rect 276 796 278 804
rect 234 795 278 796
rect 234 794 246 795
rect 266 794 278 795
rect 394 805 406 806
rect 522 805 534 806
rect 394 804 534 805
rect 394 796 396 804
rect 404 796 524 804
rect 532 796 534 804
rect 394 795 534 796
rect 394 794 406 795
rect 522 794 534 795
rect 666 805 678 806
rect 778 805 790 806
rect 666 804 790 805
rect 666 796 668 804
rect 676 796 780 804
rect 788 796 790 804
rect 666 795 790 796
rect 666 794 678 795
rect 778 794 790 795
rect 842 805 854 806
rect 1034 805 1046 806
rect 842 804 1046 805
rect 842 796 844 804
rect 852 796 1036 804
rect 1044 796 1046 804
rect 842 795 1046 796
rect 842 794 854 795
rect 1034 794 1046 795
rect 1434 805 1446 806
rect 1658 805 1670 806
rect 2122 805 2134 806
rect 1434 804 2134 805
rect 1434 796 1436 804
rect 1444 796 1660 804
rect 1668 796 2124 804
rect 2132 796 2134 804
rect 1434 795 2134 796
rect 1434 794 1446 795
rect 1658 794 1670 795
rect 2122 794 2134 795
rect 218 765 230 766
rect 314 765 326 766
rect 378 765 390 766
rect 490 765 502 766
rect -37 764 502 765
rect -37 756 220 764
rect 228 756 316 764
rect 324 756 380 764
rect 388 756 492 764
rect 500 756 502 764
rect -37 755 502 756
rect -37 715 -27 755
rect 218 754 230 755
rect 314 754 326 755
rect 378 754 390 755
rect 490 754 502 755
rect 730 765 742 766
rect 890 765 902 766
rect 730 764 902 765
rect 730 756 732 764
rect 740 756 892 764
rect 900 756 902 764
rect 730 755 902 756
rect 730 754 742 755
rect 890 754 902 755
rect 970 765 982 766
rect 1066 765 1078 766
rect 970 764 1078 765
rect 970 756 972 764
rect 980 756 1068 764
rect 1076 756 1078 764
rect 970 755 1078 756
rect 970 754 982 755
rect 1066 754 1078 755
rect 1178 765 1190 766
rect 1450 765 1462 766
rect 1178 764 1462 765
rect 1178 756 1180 764
rect 1188 756 1452 764
rect 1460 756 1462 764
rect 1178 755 1462 756
rect 1178 754 1190 755
rect 1450 754 1462 755
rect 1482 765 1494 766
rect 1546 765 1558 766
rect 1482 764 1558 765
rect 1482 756 1484 764
rect 1492 756 1548 764
rect 1556 756 1558 764
rect 1482 755 1558 756
rect 1482 754 1494 755
rect 1546 754 1558 755
rect 1578 765 1590 766
rect 1674 765 1686 766
rect 1578 764 1686 765
rect 1578 756 1580 764
rect 1588 756 1676 764
rect 1684 756 1686 764
rect 1578 755 1686 756
rect 1578 754 1590 755
rect 1674 754 1686 755
rect 1738 765 1750 766
rect 1930 765 1942 766
rect 1738 764 1942 765
rect 1738 756 1740 764
rect 1748 756 1932 764
rect 1940 756 1942 764
rect 1738 755 1942 756
rect 1738 754 1750 755
rect 1930 754 1942 755
rect 1962 765 1974 766
rect 2154 765 2166 766
rect 1962 764 2166 765
rect 1962 756 1964 764
rect 1972 756 2156 764
rect 2164 756 2166 764
rect 1962 755 2166 756
rect 1962 754 1974 755
rect 2154 754 2166 755
rect 282 725 294 726
rect 330 725 342 726
rect 282 724 342 725
rect 282 716 284 724
rect 292 716 332 724
rect 340 716 342 724
rect 282 715 342 716
rect 282 714 294 715
rect 330 714 342 715
rect 890 725 902 726
rect 922 725 934 726
rect 890 724 934 725
rect 890 716 892 724
rect 900 716 924 724
rect 932 716 934 724
rect 890 715 934 716
rect 890 714 902 715
rect 922 714 934 715
rect 1146 725 1158 726
rect 1242 725 1254 726
rect 1146 724 1254 725
rect 1146 716 1148 724
rect 1156 716 1244 724
rect 1252 716 1254 724
rect 1146 715 1254 716
rect 1146 714 1158 715
rect 1242 714 1254 715
rect 1306 725 1318 726
rect 1338 725 1350 726
rect 1306 724 1350 725
rect 1306 716 1308 724
rect 1316 716 1340 724
rect 1348 716 1350 724
rect 1306 715 1350 716
rect 1306 714 1318 715
rect 1338 714 1350 715
rect 1386 725 1398 726
rect 1482 725 1494 726
rect 1386 724 1494 725
rect 1386 716 1388 724
rect 1396 716 1484 724
rect 1492 716 1494 724
rect 1386 715 1494 716
rect 1386 714 1398 715
rect 1482 714 1494 715
rect 1514 725 1526 726
rect 1802 725 1814 726
rect 1866 725 1878 726
rect 1514 724 1878 725
rect 1514 716 1516 724
rect 1524 716 1804 724
rect 1812 716 1868 724
rect 1876 716 1878 724
rect 1514 715 1878 716
rect 1514 714 1526 715
rect 1802 714 1814 715
rect 1866 714 1878 715
rect 74 704 86 706
rect 74 696 76 704
rect 84 696 86 704
rect 74 694 86 696
rect 106 704 118 706
rect 106 696 108 704
rect 116 696 118 704
rect 106 694 118 696
rect 490 704 502 706
rect 490 696 492 704
rect 500 696 502 704
rect 490 694 502 696
rect 1130 704 1142 706
rect 1130 696 1132 704
rect 1140 696 1142 704
rect 1130 694 1142 696
rect 10 685 22 686
rect 42 685 54 686
rect 10 684 54 685
rect 10 676 12 684
rect 20 676 44 684
rect 52 676 54 684
rect 10 675 54 676
rect 10 674 22 675
rect 42 674 54 675
rect 75 645 85 694
rect 107 685 117 694
rect 218 685 230 686
rect 298 685 310 686
rect 107 675 149 685
rect 106 645 118 646
rect 75 644 118 645
rect 75 636 108 644
rect 116 636 118 644
rect 75 635 118 636
rect 139 645 149 675
rect 218 684 310 685
rect 218 676 220 684
rect 228 676 300 684
rect 308 676 310 684
rect 218 675 310 676
rect 218 674 230 675
rect 298 674 310 675
rect 330 685 342 686
rect 362 685 374 686
rect 330 684 374 685
rect 330 676 332 684
rect 340 676 364 684
rect 372 676 374 684
rect 330 675 374 676
rect 491 685 501 694
rect 650 685 662 686
rect 682 685 694 686
rect 491 684 694 685
rect 491 676 652 684
rect 660 676 684 684
rect 692 676 694 684
rect 491 675 694 676
rect 330 674 342 675
rect 362 674 374 675
rect 650 674 662 675
rect 682 674 694 675
rect 826 685 838 686
rect 858 685 870 686
rect 826 684 870 685
rect 826 676 828 684
rect 836 676 860 684
rect 868 676 870 684
rect 826 675 870 676
rect 826 674 838 675
rect 858 674 870 675
rect 906 685 918 686
rect 1018 685 1030 686
rect 906 684 1030 685
rect 906 676 908 684
rect 916 676 1020 684
rect 1028 676 1030 684
rect 906 675 1030 676
rect 906 674 918 675
rect 1018 674 1030 675
rect 1066 685 1078 686
rect 1098 685 1110 686
rect 1066 684 1110 685
rect 1066 676 1068 684
rect 1076 676 1100 684
rect 1108 676 1110 684
rect 1066 675 1110 676
rect 1131 685 1141 694
rect 1322 685 1334 686
rect 1434 685 1446 686
rect 1131 684 1446 685
rect 1131 676 1324 684
rect 1332 676 1436 684
rect 1444 676 1446 684
rect 1131 675 1446 676
rect 1066 674 1078 675
rect 1098 674 1110 675
rect 1322 674 1334 675
rect 1434 674 1446 675
rect 1674 685 1686 686
rect 1786 685 1798 686
rect 2042 685 2054 686
rect 1674 684 1717 685
rect 1674 676 1676 684
rect 1684 676 1717 684
rect 1674 675 1717 676
rect 1674 674 1686 675
rect 1707 646 1717 675
rect 1786 684 2054 685
rect 1786 676 1788 684
rect 1796 676 2044 684
rect 2052 676 2054 684
rect 1786 675 2054 676
rect 1786 674 1798 675
rect 2042 674 2054 675
rect 282 645 294 646
rect 139 644 294 645
rect 139 636 284 644
rect 292 636 294 644
rect 139 635 294 636
rect 106 634 118 635
rect 282 634 294 635
rect 314 645 326 646
rect 346 645 358 646
rect 314 644 358 645
rect 314 636 316 644
rect 324 636 348 644
rect 356 636 358 644
rect 314 635 358 636
rect 314 634 326 635
rect 346 634 358 635
rect 442 645 454 646
rect 570 645 582 646
rect 442 644 582 645
rect 442 636 444 644
rect 452 636 572 644
rect 580 636 582 644
rect 442 635 582 636
rect 442 634 454 635
rect 570 634 582 635
rect 746 645 758 646
rect 794 645 806 646
rect 746 644 806 645
rect 746 636 748 644
rect 756 636 796 644
rect 804 636 806 644
rect 746 635 806 636
rect 746 634 758 635
rect 794 634 806 635
rect 970 645 982 646
rect 1018 645 1030 646
rect 970 644 1030 645
rect 970 636 972 644
rect 980 636 1020 644
rect 1028 636 1030 644
rect 970 635 1030 636
rect 970 634 982 635
rect 1018 634 1030 635
rect 1258 645 1270 646
rect 1450 645 1462 646
rect 1258 644 1462 645
rect 1258 636 1260 644
rect 1268 636 1452 644
rect 1460 636 1462 644
rect 1258 635 1462 636
rect 1258 634 1270 635
rect 1450 634 1462 635
rect 1498 645 1510 646
rect 1610 645 1622 646
rect 1498 644 1622 645
rect 1498 636 1500 644
rect 1508 636 1612 644
rect 1620 636 1622 644
rect 1498 635 1622 636
rect 1498 634 1510 635
rect 1610 634 1622 635
rect 1642 645 1654 646
rect 1674 645 1686 646
rect 1642 644 1686 645
rect 1642 636 1644 644
rect 1652 636 1676 644
rect 1684 636 1686 644
rect 1642 635 1686 636
rect 1642 634 1654 635
rect 1674 634 1686 635
rect 1706 644 1718 646
rect 1706 636 1708 644
rect 1716 636 1718 644
rect 1706 634 1718 636
rect 1770 645 1782 646
rect 1818 645 1830 646
rect 1770 644 1830 645
rect 1770 636 1772 644
rect 1780 636 1820 644
rect 1828 636 1830 644
rect 1770 635 1830 636
rect 1770 634 1782 635
rect 1818 634 1830 635
rect 1866 645 1878 646
rect 1962 645 1974 646
rect 1866 644 1974 645
rect 1866 636 1868 644
rect 1876 636 1964 644
rect 1972 636 1974 644
rect 1866 635 1974 636
rect 1866 634 1878 635
rect 1962 634 1974 635
rect 10 605 22 606
rect -37 604 22 605
rect -37 596 12 604
rect 20 596 22 604
rect -37 595 22 596
rect -37 555 -27 595
rect 10 594 22 595
rect 106 605 118 606
rect 138 605 150 606
rect 106 604 150 605
rect 106 596 108 604
rect 116 596 140 604
rect 148 596 150 604
rect 106 595 150 596
rect 106 594 118 595
rect 138 594 150 595
rect 170 605 182 606
rect 234 605 246 606
rect 170 604 246 605
rect 170 596 172 604
rect 180 596 236 604
rect 244 596 246 604
rect 170 595 246 596
rect 170 594 182 595
rect 234 594 246 595
rect 314 605 326 606
rect 346 605 358 606
rect 314 604 358 605
rect 314 596 316 604
rect 324 596 348 604
rect 356 596 358 604
rect 314 595 358 596
rect 314 594 326 595
rect 346 594 358 595
rect 426 605 438 606
rect 538 605 550 606
rect 426 604 550 605
rect 426 596 428 604
rect 436 596 540 604
rect 548 596 550 604
rect 426 595 550 596
rect 426 594 438 595
rect 538 594 550 595
rect 890 605 902 606
rect 1082 605 1094 606
rect 1194 605 1206 606
rect 1594 605 1606 606
rect 890 604 1606 605
rect 890 596 892 604
rect 900 596 1084 604
rect 1092 596 1196 604
rect 1204 596 1596 604
rect 1604 596 1606 604
rect 890 595 1606 596
rect 890 594 902 595
rect 1082 594 1094 595
rect 1194 594 1206 595
rect 1594 594 1606 595
rect 1674 605 1686 606
rect 1786 605 1798 606
rect 1674 604 1798 605
rect 1674 596 1676 604
rect 1684 596 1788 604
rect 1796 596 1798 604
rect 1674 595 1798 596
rect 1674 594 1686 595
rect 1786 594 1798 595
rect 1818 605 1830 606
rect 1978 605 1990 606
rect 1818 604 1990 605
rect 1818 596 1820 604
rect 1828 596 1980 604
rect 1988 596 1990 604
rect 1818 595 1990 596
rect 1818 594 1830 595
rect 1978 594 1990 595
rect 2026 605 2038 606
rect 2122 605 2134 606
rect 2026 604 2134 605
rect 2026 596 2028 604
rect 2036 596 2124 604
rect 2132 596 2134 604
rect 2026 595 2134 596
rect 2026 594 2038 595
rect 2122 594 2134 595
rect 170 584 182 586
rect 170 576 172 584
rect 180 576 182 584
rect 170 574 182 576
rect 171 565 181 574
rect 139 555 181 565
rect 234 565 246 566
rect 266 565 278 566
rect 234 564 278 565
rect 234 556 236 564
rect 244 556 268 564
rect 276 556 278 564
rect 234 555 278 556
rect 26 525 38 526
rect 139 525 149 555
rect 234 554 246 555
rect 266 554 278 555
rect 298 565 310 566
rect 330 565 342 566
rect 298 564 342 565
rect 298 556 300 564
rect 308 556 332 564
rect 340 556 342 564
rect 298 555 342 556
rect 298 554 310 555
rect 330 554 342 555
rect 714 565 726 566
rect 746 565 758 566
rect 714 564 758 565
rect 714 556 716 564
rect 724 556 748 564
rect 756 556 758 564
rect 714 555 758 556
rect 714 554 726 555
rect 746 554 758 555
rect 1066 565 1078 566
rect 1194 565 1206 566
rect 1066 564 1206 565
rect 1066 556 1068 564
rect 1076 556 1196 564
rect 1204 556 1206 564
rect 1066 555 1206 556
rect 1066 554 1078 555
rect 1194 554 1206 555
rect 1466 565 1478 566
rect 1706 565 1718 566
rect 1466 564 1718 565
rect 1466 556 1468 564
rect 1476 556 1708 564
rect 1716 556 1718 564
rect 1466 555 1718 556
rect 1466 554 1478 555
rect 1706 554 1718 555
rect 1978 565 1990 566
rect 2058 565 2070 566
rect 1978 564 2070 565
rect 1978 556 1980 564
rect 1988 556 2060 564
rect 2068 556 2070 564
rect 1978 555 2070 556
rect 1978 554 1990 555
rect 2058 554 2070 555
rect -37 485 -27 525
rect 26 524 149 525
rect 26 516 28 524
rect 36 516 149 524
rect 26 515 149 516
rect 234 525 246 526
rect 282 525 294 526
rect 234 524 294 525
rect 234 516 236 524
rect 244 516 284 524
rect 292 516 294 524
rect 234 515 294 516
rect 26 514 38 515
rect 234 514 246 515
rect 282 514 294 515
rect 618 525 630 526
rect 730 525 742 526
rect 842 525 854 526
rect 618 524 854 525
rect 618 516 620 524
rect 628 516 732 524
rect 740 516 844 524
rect 852 516 854 524
rect 618 515 854 516
rect 618 514 630 515
rect 730 514 742 515
rect 842 514 854 515
rect 1130 525 1142 526
rect 1402 525 1414 526
rect 1130 524 1414 525
rect 1130 516 1132 524
rect 1140 516 1404 524
rect 1412 516 1414 524
rect 1130 515 1414 516
rect 1130 514 1142 515
rect 1402 514 1414 515
rect 1562 525 1574 526
rect 1882 525 1894 526
rect 1562 524 1894 525
rect 1562 516 1564 524
rect 1572 516 1884 524
rect 1892 516 1894 524
rect 1562 515 1894 516
rect 1562 514 1574 515
rect 1882 514 1894 515
rect 2042 525 2054 526
rect 2106 525 2118 526
rect 2042 524 2118 525
rect 2042 516 2044 524
rect 2052 516 2108 524
rect 2116 516 2118 524
rect 2042 515 2118 516
rect 2042 514 2054 515
rect 2106 514 2118 515
rect 26 485 38 486
rect -37 484 38 485
rect -37 476 28 484
rect 36 476 38 484
rect -37 475 38 476
rect 26 474 38 475
rect 122 485 134 486
rect 250 485 262 486
rect 122 484 262 485
rect 122 476 124 484
rect 132 476 252 484
rect 260 476 262 484
rect 122 475 262 476
rect 122 474 134 475
rect 250 474 262 475
rect 298 485 310 486
rect 330 485 342 486
rect 298 484 342 485
rect 298 476 300 484
rect 308 476 332 484
rect 340 476 342 484
rect 298 475 342 476
rect 298 474 310 475
rect 330 474 342 475
rect 490 485 502 486
rect 570 485 582 486
rect 490 484 582 485
rect 490 476 492 484
rect 500 476 572 484
rect 580 476 582 484
rect 490 475 582 476
rect 490 474 502 475
rect 570 474 582 475
rect 826 485 838 486
rect 954 485 966 486
rect 826 484 966 485
rect 826 476 828 484
rect 836 476 956 484
rect 964 476 966 484
rect 826 475 966 476
rect 826 474 838 475
rect 954 474 966 475
rect 986 485 998 486
rect 1018 485 1030 486
rect 986 484 1030 485
rect 986 476 988 484
rect 996 476 1020 484
rect 1028 476 1030 484
rect 986 475 1030 476
rect 986 474 998 475
rect 1018 474 1030 475
rect 1162 485 1174 486
rect 1210 485 1222 486
rect 1162 484 1222 485
rect 1162 476 1164 484
rect 1172 476 1212 484
rect 1220 476 1222 484
rect 1162 475 1222 476
rect 1162 474 1174 475
rect 1210 474 1222 475
rect 1242 485 1254 486
rect 1370 485 1382 486
rect 1242 484 1382 485
rect 1242 476 1244 484
rect 1252 476 1372 484
rect 1380 476 1382 484
rect 1242 475 1382 476
rect 1242 474 1254 475
rect 1370 474 1382 475
rect 1466 485 1478 486
rect 1514 485 1526 486
rect 1466 484 1526 485
rect 1466 476 1468 484
rect 1476 476 1516 484
rect 1524 476 1526 484
rect 1466 475 1526 476
rect 1466 474 1478 475
rect 1514 474 1526 475
rect 1626 485 1638 486
rect 1722 485 1734 486
rect 1626 484 1734 485
rect 1626 476 1628 484
rect 1636 476 1724 484
rect 1732 476 1734 484
rect 1626 475 1734 476
rect 1626 474 1638 475
rect 1722 474 1734 475
rect 1914 485 1926 486
rect 1994 485 2006 486
rect 1914 484 2006 485
rect 1914 476 1916 484
rect 1924 476 1996 484
rect 2004 476 2006 484
rect 1914 475 2006 476
rect 1914 474 1926 475
rect 1994 474 2006 475
rect 1674 464 1686 466
rect 1674 456 1676 464
rect 1684 456 1686 464
rect 1674 454 1686 456
rect 138 445 150 446
rect 266 445 278 446
rect 138 444 278 445
rect 138 436 140 444
rect 148 436 268 444
rect 276 436 278 444
rect 138 435 278 436
rect 138 434 150 435
rect 266 434 278 435
rect 314 445 326 446
rect 346 445 358 446
rect 314 444 358 445
rect 314 436 316 444
rect 324 436 348 444
rect 356 436 358 444
rect 314 435 358 436
rect 314 434 326 435
rect 346 434 358 435
rect 378 445 390 446
rect 458 445 470 446
rect 378 444 470 445
rect 378 436 380 444
rect 388 436 460 444
rect 468 436 470 444
rect 378 435 470 436
rect 378 434 390 435
rect 458 434 470 435
rect 714 445 726 446
rect 1050 445 1062 446
rect 1082 445 1094 446
rect 714 444 1094 445
rect 714 436 716 444
rect 724 436 1052 444
rect 1060 436 1084 444
rect 1092 436 1094 444
rect 714 435 1094 436
rect 714 434 726 435
rect 1050 434 1062 435
rect 1082 434 1094 435
rect 1114 445 1126 446
rect 1194 445 1206 446
rect 1114 444 1206 445
rect 1114 436 1116 444
rect 1124 436 1196 444
rect 1204 436 1206 444
rect 1114 435 1206 436
rect 1114 434 1126 435
rect 1194 434 1206 435
rect 1370 445 1382 446
rect 1562 445 1574 446
rect 1370 444 1574 445
rect 1370 436 1372 444
rect 1380 436 1564 444
rect 1572 436 1574 444
rect 1370 435 1574 436
rect 1370 434 1382 435
rect 1562 434 1574 435
rect 1594 445 1606 446
rect 1675 445 1685 454
rect 1594 444 1685 445
rect 1594 436 1596 444
rect 1604 436 1685 444
rect 1594 435 1685 436
rect 1722 445 1734 446
rect 1802 445 1814 446
rect 1722 444 1814 445
rect 1722 436 1724 444
rect 1732 436 1804 444
rect 1812 436 1814 444
rect 1722 435 1814 436
rect 1594 434 1606 435
rect 1722 434 1734 435
rect 1802 434 1814 435
rect 1866 445 1878 446
rect 1930 445 1942 446
rect 1866 444 1942 445
rect 1866 436 1868 444
rect 1876 436 1932 444
rect 1940 436 1942 444
rect 1866 435 1942 436
rect 1866 434 1878 435
rect 1930 434 1942 435
rect 10 405 22 406
rect 58 405 70 406
rect 10 404 70 405
rect 10 396 12 404
rect 20 396 60 404
rect 68 396 70 404
rect 10 395 70 396
rect 10 394 22 395
rect 58 394 70 395
rect 186 405 198 406
rect 410 405 422 406
rect 442 405 454 406
rect 186 404 454 405
rect 186 396 188 404
rect 196 396 412 404
rect 420 396 444 404
rect 452 396 454 404
rect 186 395 454 396
rect 186 394 198 395
rect 410 394 422 395
rect 442 394 454 395
rect 554 405 566 406
rect 586 405 598 406
rect 554 404 598 405
rect 554 396 556 404
rect 564 396 588 404
rect 596 396 598 404
rect 554 395 598 396
rect 554 394 566 395
rect 586 394 598 395
rect 778 405 790 406
rect 906 405 918 406
rect 778 404 918 405
rect 778 396 780 404
rect 788 396 908 404
rect 916 396 918 404
rect 778 395 918 396
rect 778 394 790 395
rect 906 394 918 395
rect 1018 405 1030 406
rect 1082 405 1094 406
rect 1018 404 1094 405
rect 1018 396 1020 404
rect 1028 396 1084 404
rect 1092 396 1094 404
rect 1018 395 1094 396
rect 1018 394 1030 395
rect 1082 394 1094 395
rect 1306 405 1318 406
rect 1418 405 1430 406
rect 1546 405 1558 406
rect 1306 404 1558 405
rect 1306 396 1308 404
rect 1316 396 1420 404
rect 1428 396 1548 404
rect 1556 396 1558 404
rect 1306 395 1558 396
rect 1306 394 1318 395
rect 1418 394 1430 395
rect 1546 394 1558 395
rect 1610 405 1622 406
rect 1674 405 1686 406
rect 1610 404 1686 405
rect 1610 396 1612 404
rect 1620 396 1676 404
rect 1684 396 1686 404
rect 1610 395 1686 396
rect 1610 394 1622 395
rect 1674 394 1686 395
rect 1706 405 1718 406
rect 1898 405 1910 406
rect 1706 404 1910 405
rect 1706 396 1708 404
rect 1716 396 1900 404
rect 1908 396 1910 404
rect 1706 395 1910 396
rect 1706 394 1718 395
rect 1898 394 1910 395
rect 1930 405 1942 406
rect 1978 405 1990 406
rect 1930 404 1990 405
rect 1930 396 1932 404
rect 1940 396 1980 404
rect 1988 396 1990 404
rect 1930 395 1990 396
rect 1930 394 1942 395
rect 1978 394 1990 395
rect 58 365 70 366
rect 218 365 230 366
rect 58 364 230 365
rect 58 356 60 364
rect 68 356 220 364
rect 228 356 230 364
rect 58 355 230 356
rect 58 354 70 355
rect 218 354 230 355
rect 298 365 310 366
rect 362 365 374 366
rect 298 364 374 365
rect 298 356 300 364
rect 308 356 364 364
rect 372 356 374 364
rect 298 355 374 356
rect 298 354 310 355
rect 362 354 374 355
rect 410 365 422 366
rect 570 365 582 366
rect 602 365 614 366
rect 410 364 614 365
rect 410 356 412 364
rect 420 356 572 364
rect 580 356 604 364
rect 612 356 614 364
rect 410 355 614 356
rect 410 354 422 355
rect 570 354 582 355
rect 602 354 614 355
rect 1002 365 1014 366
rect 1226 365 1238 366
rect 1002 364 1238 365
rect 1002 356 1004 364
rect 1012 356 1228 364
rect 1236 356 1238 364
rect 1002 355 1238 356
rect 1002 354 1014 355
rect 1226 354 1238 355
rect 1258 365 1270 366
rect 1290 365 1302 366
rect 1258 364 1302 365
rect 1258 356 1260 364
rect 1268 356 1292 364
rect 1300 356 1302 364
rect 1258 355 1302 356
rect 1258 354 1270 355
rect 1290 354 1302 355
rect 1402 365 1414 366
rect 1642 365 1654 366
rect 1402 364 1654 365
rect 1402 356 1404 364
rect 1412 356 1644 364
rect 1652 356 1654 364
rect 1402 355 1654 356
rect 1402 354 1414 355
rect 1642 354 1654 355
rect 1786 365 1798 366
rect 1834 365 1846 366
rect 1930 365 1942 366
rect 1786 364 1846 365
rect 1786 356 1788 364
rect 1796 356 1836 364
rect 1844 356 1846 364
rect 1786 355 1846 356
rect 1786 354 1798 355
rect 1834 354 1846 355
rect 1867 364 1942 365
rect 1867 356 1932 364
rect 1940 356 1942 364
rect 1867 355 1942 356
rect 74 325 86 326
rect 106 325 118 326
rect 74 324 118 325
rect 74 316 76 324
rect 84 316 108 324
rect 116 316 118 324
rect 74 315 118 316
rect 74 314 86 315
rect 106 314 118 315
rect 218 325 230 326
rect 250 325 262 326
rect 218 324 262 325
rect 218 316 220 324
rect 228 316 252 324
rect 260 316 262 324
rect 218 315 262 316
rect 218 314 230 315
rect 250 314 262 315
rect 586 325 598 326
rect 698 325 710 326
rect 586 324 710 325
rect 586 316 588 324
rect 596 316 700 324
rect 708 316 710 324
rect 586 315 710 316
rect 586 314 598 315
rect 698 314 710 315
rect 746 325 758 326
rect 810 325 822 326
rect 842 325 854 326
rect 1104 325 1126 326
rect 746 324 854 325
rect 746 316 748 324
rect 756 316 812 324
rect 820 316 844 324
rect 852 316 854 324
rect 746 315 854 316
rect 746 314 758 315
rect 810 314 822 315
rect 842 314 854 315
rect 1099 324 1126 325
rect 1099 316 1116 324
rect 1124 316 1126 324
rect 1099 314 1126 316
rect 1226 325 1238 326
rect 1322 325 1334 326
rect 1226 324 1334 325
rect 1226 316 1228 324
rect 1236 316 1324 324
rect 1332 316 1334 324
rect 1226 315 1334 316
rect 1226 314 1238 315
rect 1322 314 1334 315
rect 1466 325 1478 326
rect 1546 325 1558 326
rect 1466 324 1558 325
rect 1466 316 1468 324
rect 1476 316 1548 324
rect 1556 316 1558 324
rect 1466 315 1558 316
rect 1466 314 1478 315
rect 1546 314 1558 315
rect 1658 325 1670 326
rect 1690 325 1702 326
rect 1658 324 1702 325
rect 1658 316 1660 324
rect 1668 316 1692 324
rect 1700 316 1702 324
rect 1658 315 1702 316
rect 1658 314 1670 315
rect 1690 314 1702 315
rect 1786 325 1798 326
rect 1867 325 1877 355
rect 1930 354 1942 355
rect 2090 365 2102 366
rect 2154 365 2166 366
rect 2090 364 2166 365
rect 2090 356 2092 364
rect 2100 356 2156 364
rect 2164 356 2166 364
rect 2090 355 2166 356
rect 2090 354 2102 355
rect 2154 354 2166 355
rect 1786 324 1877 325
rect 1786 316 1788 324
rect 1796 316 1877 324
rect 1786 315 1877 316
rect 2026 325 2038 326
rect 2074 325 2086 326
rect 2026 324 2086 325
rect 2026 316 2028 324
rect 2036 316 2076 324
rect 2084 316 2086 324
rect 2026 315 2086 316
rect 1786 314 1798 315
rect 2026 314 2038 315
rect 2074 314 2086 315
rect 2106 325 2118 326
rect 2203 325 2213 345
rect 2106 324 2213 325
rect 2106 316 2108 324
rect 2116 316 2213 324
rect 2106 315 2213 316
rect 2106 314 2118 315
rect 10 285 22 286
rect 138 285 150 286
rect 10 284 150 285
rect 10 276 12 284
rect 20 276 140 284
rect 148 276 150 284
rect 10 275 150 276
rect 10 274 22 275
rect 138 274 150 275
rect 234 285 246 286
rect 346 285 358 286
rect 714 285 726 286
rect 826 285 838 286
rect 1099 285 1109 314
rect 1290 304 1302 306
rect 1290 296 1292 304
rect 1300 296 1302 304
rect 1290 294 1302 296
rect 1770 304 1782 306
rect 1770 296 1772 304
rect 1780 296 1782 304
rect 1770 294 1782 296
rect 1291 285 1301 294
rect 234 284 358 285
rect 234 276 236 284
rect 244 276 348 284
rect 356 276 358 284
rect 234 275 358 276
rect 234 274 246 275
rect 346 274 358 275
rect 587 284 1109 285
rect 587 276 716 284
rect 724 276 828 284
rect 836 276 1109 284
rect 587 275 1109 276
rect 1227 275 1301 285
rect 1546 285 1558 286
rect 1658 285 1670 286
rect 1546 284 1670 285
rect 1546 276 1548 284
rect 1556 276 1660 284
rect 1668 276 1670 284
rect 1546 275 1670 276
rect 587 266 597 275
rect 714 274 726 275
rect 826 274 838 275
rect 586 264 598 266
rect 586 256 588 264
rect 596 256 598 264
rect 586 254 598 256
rect 362 245 374 246
rect 490 245 502 246
rect 362 244 502 245
rect 362 236 364 244
rect 372 236 492 244
rect 500 236 502 244
rect 362 235 502 236
rect 362 234 374 235
rect 490 234 502 235
rect 714 245 726 246
rect 794 245 806 246
rect 714 244 806 245
rect 714 236 716 244
rect 724 236 796 244
rect 804 236 806 244
rect 714 235 806 236
rect 714 234 726 235
rect 794 234 806 235
rect 874 245 886 246
rect 970 245 982 246
rect 874 244 982 245
rect 874 236 876 244
rect 884 236 972 244
rect 980 236 982 244
rect 874 235 982 236
rect 874 234 886 235
rect 970 234 982 235
rect 1002 245 1014 246
rect 1034 245 1046 246
rect 1002 244 1046 245
rect 1002 236 1004 244
rect 1012 236 1036 244
rect 1044 236 1046 244
rect 1002 235 1046 236
rect 1002 234 1014 235
rect 1034 234 1046 235
rect 1146 245 1158 246
rect 1227 245 1237 275
rect 1546 274 1558 275
rect 1658 274 1670 275
rect 1771 246 1781 294
rect 1850 285 1862 286
rect 1914 285 1926 286
rect 1850 284 1926 285
rect 1850 276 1852 284
rect 1860 276 1916 284
rect 1924 276 1926 284
rect 1850 275 1926 276
rect 1850 274 1862 275
rect 1914 274 1926 275
rect 1946 285 1958 286
rect 2058 285 2070 286
rect 1946 284 2070 285
rect 1946 276 1948 284
rect 1956 276 2060 284
rect 2068 276 2070 284
rect 1946 275 2070 276
rect 1946 274 1958 275
rect 2058 274 2070 275
rect 2154 285 2166 286
rect 2203 285 2213 305
rect 2154 284 2213 285
rect 2154 276 2156 284
rect 2164 276 2213 284
rect 2154 275 2213 276
rect 2154 274 2166 275
rect 1146 244 1237 245
rect 1146 236 1148 244
rect 1156 236 1237 244
rect 1146 235 1237 236
rect 1258 245 1270 246
rect 1370 245 1382 246
rect 1258 244 1382 245
rect 1258 236 1260 244
rect 1268 236 1372 244
rect 1380 236 1382 244
rect 1258 235 1382 236
rect 1146 234 1158 235
rect 1258 234 1270 235
rect 1370 234 1382 235
rect 1514 245 1526 246
rect 1594 245 1606 246
rect 1514 244 1606 245
rect 1514 236 1516 244
rect 1524 236 1596 244
rect 1604 236 1606 244
rect 1514 235 1606 236
rect 1514 234 1526 235
rect 1594 234 1606 235
rect 1642 245 1654 246
rect 1674 245 1686 246
rect 1642 244 1686 245
rect 1642 236 1644 244
rect 1652 236 1676 244
rect 1684 236 1686 244
rect 1642 235 1686 236
rect 1642 234 1654 235
rect 1674 234 1686 235
rect 1770 244 1782 246
rect 1770 236 1772 244
rect 1780 236 1782 244
rect 1770 234 1782 236
rect 1882 245 1894 246
rect 1946 245 1958 246
rect 1882 244 1958 245
rect 1882 236 1884 244
rect 1892 236 1948 244
rect 1956 236 1958 244
rect 1882 235 1958 236
rect 1882 234 1894 235
rect 1946 234 1958 235
rect 106 205 118 206
rect 202 205 214 206
rect 106 204 214 205
rect 106 196 108 204
rect 116 196 204 204
rect 212 196 214 204
rect 106 195 214 196
rect 106 194 118 195
rect 202 194 214 195
rect 730 205 742 206
rect 1178 205 1190 206
rect 730 204 1190 205
rect 730 196 732 204
rect 740 196 1180 204
rect 1188 196 1190 204
rect 730 195 1190 196
rect 730 194 742 195
rect 1178 194 1190 195
rect 1418 205 1430 206
rect 1546 205 1558 206
rect 1418 204 1558 205
rect 1418 196 1420 204
rect 1428 196 1548 204
rect 1556 196 1558 204
rect 1418 195 1558 196
rect 1418 194 1430 195
rect 1546 194 1558 195
rect 1690 205 1702 206
rect 1722 205 1734 206
rect 1690 204 1734 205
rect 1690 196 1692 204
rect 1700 196 1724 204
rect 1732 196 1734 204
rect 1690 195 1734 196
rect 1690 194 1702 195
rect 1722 194 1734 195
rect 1754 205 1766 206
rect 1802 205 1814 206
rect 1754 204 1814 205
rect 1754 196 1756 204
rect 1764 196 1804 204
rect 1812 196 1814 204
rect 1754 195 1814 196
rect 1754 194 1766 195
rect 1802 194 1814 195
rect 1962 205 1974 206
rect 2026 205 2038 206
rect 1962 204 2038 205
rect 1962 196 1964 204
rect 1972 196 2028 204
rect 2036 196 2038 204
rect 1962 195 2038 196
rect 1962 194 1974 195
rect 2026 194 2038 195
rect 218 165 230 166
rect 346 165 358 166
rect 218 164 358 165
rect 218 156 220 164
rect 228 156 348 164
rect 356 156 358 164
rect 218 155 358 156
rect 218 154 230 155
rect 346 154 358 155
rect 490 165 502 166
rect 602 165 614 166
rect 778 165 790 166
rect 1114 165 1126 166
rect 490 164 614 165
rect 490 156 492 164
rect 500 156 604 164
rect 612 156 614 164
rect 490 155 614 156
rect 490 154 502 155
rect 602 154 614 155
rect 651 164 790 165
rect 651 156 780 164
rect 788 156 790 164
rect 651 155 790 156
rect 10 125 22 126
rect 122 125 134 126
rect 186 125 198 126
rect 10 124 198 125
rect 10 116 12 124
rect 20 116 124 124
rect 132 116 188 124
rect 196 116 198 124
rect 10 115 198 116
rect 10 114 22 115
rect 122 114 134 115
rect 186 114 198 115
rect 250 125 262 126
rect 314 125 326 126
rect 250 124 326 125
rect 250 116 252 124
rect 260 116 316 124
rect 324 116 326 124
rect 250 115 326 116
rect 250 114 262 115
rect 314 114 326 115
rect 362 125 374 126
rect 474 125 486 126
rect 362 124 486 125
rect 362 116 364 124
rect 372 116 476 124
rect 484 116 486 124
rect 362 115 486 116
rect 362 114 374 115
rect 474 114 486 115
rect 602 125 614 126
rect 651 125 661 155
rect 778 154 790 155
rect 1035 164 1126 165
rect 1035 156 1116 164
rect 1124 156 1126 164
rect 1035 155 1126 156
rect 602 124 661 125
rect 602 116 604 124
rect 612 116 661 124
rect 602 115 661 116
rect 698 125 710 126
rect 762 125 774 126
rect 826 125 838 126
rect 698 124 838 125
rect 698 116 700 124
rect 708 116 764 124
rect 772 116 828 124
rect 836 116 838 124
rect 698 115 838 116
rect 602 114 614 115
rect 698 114 710 115
rect 762 114 774 115
rect 826 114 838 115
rect 906 125 918 126
rect 1035 125 1045 155
rect 1114 154 1126 155
rect 1146 165 1158 166
rect 1322 165 1334 166
rect 1146 164 1334 165
rect 1146 156 1148 164
rect 1156 156 1324 164
rect 1332 156 1334 164
rect 1146 155 1334 156
rect 1146 154 1158 155
rect 1322 154 1334 155
rect 1594 165 1606 166
rect 1706 165 1718 166
rect 1754 165 1766 166
rect 1594 164 1653 165
rect 1594 156 1596 164
rect 1604 156 1653 164
rect 1594 155 1653 156
rect 1594 154 1606 155
rect 906 124 1045 125
rect 906 116 908 124
rect 916 116 1045 124
rect 906 115 1045 116
rect 1098 125 1110 126
rect 1146 125 1158 126
rect 1098 124 1158 125
rect 1098 116 1100 124
rect 1108 116 1148 124
rect 1156 116 1158 124
rect 1098 115 1158 116
rect 906 114 918 115
rect 1098 114 1110 115
rect 1146 114 1158 115
rect 1178 125 1190 126
rect 1210 125 1222 126
rect 1178 124 1222 125
rect 1178 116 1180 124
rect 1188 116 1212 124
rect 1220 116 1222 124
rect 1178 115 1222 116
rect 1178 114 1190 115
rect 1210 114 1222 115
rect 1290 125 1302 126
rect 1530 125 1542 126
rect 1290 124 1542 125
rect 1290 116 1292 124
rect 1300 116 1532 124
rect 1540 116 1542 124
rect 1290 115 1542 116
rect 1290 114 1302 115
rect 1530 114 1542 115
rect 1562 125 1574 126
rect 1610 125 1622 126
rect 1562 124 1622 125
rect 1562 116 1564 124
rect 1572 116 1612 124
rect 1620 116 1622 124
rect 1562 115 1622 116
rect 1643 125 1653 155
rect 1706 164 1766 165
rect 1706 156 1708 164
rect 1716 156 1756 164
rect 1764 156 1766 164
rect 1706 155 1766 156
rect 1706 154 1718 155
rect 1754 154 1766 155
rect 1802 165 1814 166
rect 2122 165 2134 166
rect 1802 164 2134 165
rect 1802 156 1804 164
rect 1812 156 2124 164
rect 2132 156 2134 164
rect 1802 155 2134 156
rect 1802 154 1814 155
rect 2122 154 2134 155
rect 1690 125 1702 126
rect 1643 124 1702 125
rect 1643 116 1692 124
rect 1700 116 1702 124
rect 1643 115 1702 116
rect 1562 114 1574 115
rect 1610 114 1622 115
rect 1690 114 1702 115
rect 1738 125 1750 126
rect 1834 125 1846 126
rect 1738 124 1846 125
rect 1738 116 1740 124
rect 1748 116 1836 124
rect 1844 116 1846 124
rect 1738 115 1846 116
rect 1738 114 1750 115
rect 1834 114 1846 115
rect 1914 125 1926 126
rect 2090 125 2102 126
rect 1914 124 2102 125
rect 1914 116 1916 124
rect 1924 116 2092 124
rect 2100 116 2102 124
rect 1914 115 2102 116
rect 1914 114 1926 115
rect 2090 114 2102 115
rect 106 85 118 86
rect 218 85 230 86
rect 106 84 230 85
rect 106 76 108 84
rect 116 76 220 84
rect 228 76 230 84
rect 106 75 230 76
rect 106 74 118 75
rect 218 74 230 75
rect 298 85 310 86
rect 778 85 790 86
rect 298 84 790 85
rect 298 76 300 84
rect 308 76 780 84
rect 788 76 790 84
rect 298 75 790 76
rect 298 74 310 75
rect 778 74 790 75
rect 810 85 822 86
rect 1354 85 1366 86
rect 810 84 1366 85
rect 810 76 812 84
rect 820 76 1356 84
rect 1364 76 1366 84
rect 810 75 1366 76
rect 810 74 822 75
rect 1354 74 1366 75
rect 1386 85 1398 86
rect 1418 85 1430 86
rect 1386 84 1430 85
rect 1386 76 1388 84
rect 1396 76 1420 84
rect 1428 76 1430 84
rect 1386 75 1430 76
rect 1386 74 1398 75
rect 1418 74 1430 75
rect 1482 85 1494 86
rect 1546 85 1558 86
rect 1482 84 1558 85
rect 1482 76 1484 84
rect 1492 76 1548 84
rect 1556 76 1558 84
rect 1482 75 1558 76
rect 1482 74 1494 75
rect 1546 74 1558 75
rect 1754 85 1766 86
rect 1914 85 1926 86
rect 1754 84 1926 85
rect 1754 76 1756 84
rect 1764 76 1916 84
rect 1924 76 1926 84
rect 1754 75 1926 76
rect 1754 74 1766 75
rect 1914 74 1926 75
rect 650 45 662 46
rect 698 45 710 46
rect 650 44 710 45
rect 650 36 652 44
rect 660 36 700 44
rect 708 36 710 44
rect 650 35 710 36
rect 650 34 662 35
rect 698 34 710 35
rect 730 45 742 46
rect 794 45 806 46
rect 730 44 806 45
rect 730 36 732 44
rect 740 36 796 44
rect 804 36 806 44
rect 730 35 806 36
rect 730 34 742 35
rect 794 34 806 35
rect 826 45 838 46
rect 906 45 918 46
rect 826 44 918 45
rect 826 36 828 44
rect 836 36 908 44
rect 916 36 918 44
rect 826 35 918 36
rect 826 34 838 35
rect 906 34 918 35
rect 1002 45 1014 46
rect 1034 45 1046 46
rect 1162 45 1174 46
rect 1002 44 1046 45
rect 1002 36 1004 44
rect 1012 36 1036 44
rect 1044 36 1046 44
rect 1002 35 1046 36
rect 1002 34 1014 35
rect 1034 34 1046 35
rect 1067 44 1174 45
rect 1067 36 1164 44
rect 1172 36 1174 44
rect 1067 35 1174 36
rect 1067 26 1077 35
rect 1162 34 1174 35
rect 1242 45 1254 46
rect 1306 45 1318 46
rect 1242 44 1318 45
rect 1242 36 1244 44
rect 1252 36 1308 44
rect 1316 36 1318 44
rect 1242 35 1318 36
rect 1242 34 1254 35
rect 1306 34 1318 35
rect 1338 45 1350 46
rect 1370 45 1382 46
rect 1338 44 1382 45
rect 1338 36 1340 44
rect 1348 36 1372 44
rect 1380 36 1382 44
rect 1338 35 1382 36
rect 1338 34 1350 35
rect 1370 34 1382 35
rect 1594 45 1606 46
rect 1674 45 1686 46
rect 1594 44 1686 45
rect 1594 36 1596 44
rect 1604 36 1676 44
rect 1684 36 1686 44
rect 1594 35 1686 36
rect 1594 34 1606 35
rect 1674 34 1686 35
rect 1706 45 1718 46
rect 2026 45 2038 46
rect 1706 44 2038 45
rect 1706 36 1708 44
rect 1716 36 2028 44
rect 2036 36 2038 44
rect 1706 35 2038 36
rect 1706 34 1718 35
rect 2026 34 2038 35
rect 1066 24 1078 26
rect 1066 16 1068 24
rect 1076 16 1078 24
rect 1066 14 1078 16
use AND2X2  _104_
timestamp 1656222261
transform 1 0 8 0 -1 1410
box 0 0 64 200
use AND2X2  _103_
timestamp 1656222261
transform -1 0 136 0 -1 1410
box 0 0 64 200
use XOR2X1  _125_
timestamp 1656222261
transform -1 0 248 0 -1 1410
box 0 0 112 200
use AND2X2  _126_
timestamp 1656222261
transform 1 0 248 0 -1 1410
box 0 0 64 200
use OR2X2  _124_
timestamp 1656222261
transform 1 0 312 0 -1 1410
box 0 0 64 200
use AND2X2  _100_
timestamp 1656222261
transform -1 0 440 0 -1 1410
box 0 0 64 200
use AND2X2  _97_
timestamp 1656222261
transform 1 0 440 0 -1 1410
box 0 0 64 200
use AND2X2  _99_
timestamp 1656222261
transform 1 0 504 0 -1 1410
box 0 0 64 200
use AND2X2  _108_
timestamp 1656222261
transform 1 0 568 0 -1 1410
box 0 0 64 200
use XOR2X1  _107_
timestamp 1656222261
transform -1 0 744 0 -1 1410
box 0 0 112 200
use BUFX2  _0_
timestamp 1656222261
transform -1 0 792 0 -1 1410
box 0 0 48 200
use DFFSR  _9_
timestamp 1656222261
transform -1 0 1144 0 -1 1410
box 0 0 352 200
use XOR2X1  _24_
timestamp 1656222261
transform -1 0 1256 0 -1 1410
box 0 0 112 200
use AND2X2  _25_
timestamp 1656222261
transform -1 0 1320 0 -1 1410
box 0 0 64 200
use BUFX2  _1_
timestamp 1656222261
transform -1 0 1368 0 -1 1410
box 0 0 48 200
use DFFSR  _10_
timestamp 1656222261
transform -1 0 1720 0 -1 1410
box 0 0 352 200
use DFFSR  _11_
timestamp 1656222261
transform 1 0 1720 0 -1 1410
box 0 0 352 200
use BUFX2  _2_
timestamp 1656222261
transform 1 0 2072 0 -1 1410
box 0 0 48 200
use FILL  FILL31800x18150
timestamp 1656222261
transform -1 0 2136 0 -1 1410
box 0 0 16 200
use FILL  FILL32040x18150
timestamp 1656222261
transform -1 0 2152 0 -1 1410
box 0 0 16 200
use FILL  FILL32280x18150
timestamp 1656222261
transform -1 0 2168 0 -1 1410
box 0 0 16 200
use XOR2X1  _130_
timestamp 1656222261
transform 1 0 8 0 1 1010
box 0 0 112 200
use AND2X2  _131_
timestamp 1656222261
transform 1 0 120 0 1 1010
box 0 0 64 200
use AND2X2  _91_
timestamp 1656222261
transform -1 0 248 0 1 1010
box 0 0 64 200
use AND2X2  _95_
timestamp 1656222261
transform 1 0 248 0 1 1010
box 0 0 64 200
use AND2X2  _128_
timestamp 1656222261
transform -1 0 376 0 1 1010
box 0 0 64 200
use XOR2X1  _127_
timestamp 1656222261
transform -1 0 488 0 1 1010
box 0 0 112 200
use AND2X2  _96_
timestamp 1656222261
transform 1 0 488 0 1 1010
box 0 0 64 200
use XOR2X1  _136_
timestamp 1656222261
transform -1 0 664 0 1 1010
box 0 0 112 200
use AND2X2  _137_
timestamp 1656222261
transform 1 0 664 0 1 1010
box 0 0 64 200
use XOR2X1  _19_
timestamp 1656222261
transform -1 0 840 0 1 1010
box 0 0 112 200
use AND2X2  _20_
timestamp 1656222261
transform 1 0 840 0 1 1010
box 0 0 64 200
use OR2X2  _18_
timestamp 1656222261
transform 1 0 904 0 1 1010
box 0 0 64 200
use AND2X2  _22_
timestamp 1656222261
transform -1 0 1032 0 1 1010
box 0 0 64 200
use XOR2X1  _21_
timestamp 1656222261
transform -1 0 1144 0 1 1010
box 0 0 112 200
use AND2X2  _27_
timestamp 1656222261
transform 1 0 1144 0 1 1010
box 0 0 64 200
use OR2X2  _23_
timestamp 1656222261
transform 1 0 1208 0 1 1010
box 0 0 64 200
use XOR2X1  _26_
timestamp 1656222261
transform -1 0 1384 0 1 1010
box 0 0 112 200
use XOR2X1  _84_
timestamp 1656222261
transform -1 0 1496 0 1 1010
box 0 0 112 200
use AND2X2  _85_
timestamp 1656222261
transform 1 0 1496 0 1 1010
box 0 0 64 200
use AND2X2  _90_
timestamp 1656222261
transform 1 0 1560 0 1 1010
box 0 0 64 200
use AND2X2  _88_
timestamp 1656222261
transform 1 0 1624 0 1 1010
box 0 0 64 200
use XOR2X1  _87_
timestamp 1656222261
transform -1 0 1800 0 1 1010
box 0 0 112 200
use XOR2X1  _89_
timestamp 1656222261
transform 1 0 1800 0 1 1010
box 0 0 112 200
use XOR2X1  _57_
timestamp 1656222261
transform 1 0 1912 0 1 1010
box 0 0 112 200
use XOR2X1  _55_
timestamp 1656222261
transform -1 0 2136 0 1 1010
box 0 0 112 200
use FILL  FILL32040x15150
timestamp 1656222261
transform 1 0 2136 0 1 1010
box 0 0 16 200
use FILL  FILL32280x15150
timestamp 1656222261
transform 1 0 2152 0 1 1010
box 0 0 16 200
use XOR2X1  _132_
timestamp 1656222261
transform -1 0 120 0 -1 1010
box 0 0 112 200
use AND2X2  _133_
timestamp 1656222261
transform 1 0 120 0 -1 1010
box 0 0 64 200
use OR2X2  _129_
timestamp 1656222261
transform 1 0 184 0 -1 1010
box 0 0 64 200
use AND2X2  _101_
timestamp 1656222261
transform -1 0 312 0 -1 1010
box 0 0 64 200
use XOR2X1  _139_
timestamp 1656222261
transform -1 0 424 0 -1 1010
box 0 0 112 200
use AND2X2  _140_
timestamp 1656222261
transform 1 0 424 0 -1 1010
box 0 0 64 200
use AND2X2  _98_
timestamp 1656222261
transform 1 0 488 0 -1 1010
box 0 0 64 200
use OR2X2  _138_
timestamp 1656222261
transform -1 0 616 0 -1 1010
box 0 0 64 200
use AND2X2  _142_
timestamp 1656222261
transform -1 0 680 0 -1 1010
box 0 0 64 200
use XOR2X1  _141_
timestamp 1656222261
transform 1 0 680 0 -1 1010
box 0 0 112 200
use AND2X2  _154_
timestamp 1656222261
transform -1 0 856 0 -1 1010
box 0 0 64 200
use XOR2X1  _153_
timestamp 1656222261
transform 1 0 856 0 -1 1010
box 0 0 112 200
use DFFSR  _13_
timestamp 1656222261
transform -1 0 1320 0 -1 1010
box 0 0 352 200
use OR2X2  _59_
timestamp 1656222261
transform -1 0 1384 0 -1 1010
box 0 0 64 200
use AND2X2  _61_
timestamp 1656222261
transform -1 0 1448 0 -1 1010
box 0 0 64 200
use AND2X2  _63_
timestamp 1656222261
transform -1 0 1512 0 -1 1010
box 0 0 64 200
use BUFX2  BUFX2_insert0
timestamp 1656222261
transform -1 0 1560 0 -1 1010
box 0 0 48 200
use XOR2X1  _60_
timestamp 1656222261
transform -1 0 1672 0 -1 1010
box 0 0 112 200
use OR2X2  _86_
timestamp 1656222261
transform 1 0 1672 0 -1 1010
box 0 0 64 200
use BUFX2  BUFX2_insert2
timestamp 1656222261
transform 1 0 1736 0 -1 1010
box 0 0 48 200
use XOR2X1  _62_
timestamp 1656222261
transform -1 0 1896 0 -1 1010
box 0 0 112 200
use OR2X2  _54_
timestamp 1656222261
transform -1 0 1960 0 -1 1010
box 0 0 64 200
use AND2X2  _58_
timestamp 1656222261
transform -1 0 2024 0 -1 1010
box 0 0 64 200
use BUFX2  _8_
timestamp 1656222261
transform 1 0 2024 0 -1 1010
box 0 0 48 200
use AND2X2  _56_
timestamp 1656222261
transform -1 0 2136 0 -1 1010
box 0 0 64 200
use FILL  FILL32040x12150
timestamp 1656222261
transform -1 0 2152 0 -1 1010
box 0 0 16 200
use FILL  FILL32280x12150
timestamp 1656222261
transform -1 0 2168 0 -1 1010
box 0 0 16 200
use AND2X2  _92_
timestamp 1656222261
transform 1 0 8 0 1 610
box 0 0 64 200
use XOR2X1  _134_
timestamp 1656222261
transform -1 0 184 0 1 610
box 0 0 112 200
use AND2X2  _94_
timestamp 1656222261
transform -1 0 248 0 1 610
box 0 0 64 200
use AND2X2  _105_
timestamp 1656222261
transform -1 0 312 0 1 610
box 0 0 64 200
use AND2X2  _106_
timestamp 1656222261
transform 1 0 312 0 1 610
box 0 0 64 200
use AND2X2  _102_
timestamp 1656222261
transform 1 0 376 0 1 610
box 0 0 64 200
use XOR2X1  _110_
timestamp 1656222261
transform -1 0 552 0 1 610
box 0 0 112 200
use AND2X2  _111_
timestamp 1656222261
transform 1 0 552 0 1 610
box 0 0 64 200
use AND2X2  _113_
timestamp 1656222261
transform -1 0 680 0 1 610
box 0 0 64 200
use XOR2X1  _112_
timestamp 1656222261
transform -1 0 792 0 1 610
box 0 0 112 200
use OR2X2  _64_
timestamp 1656222261
transform -1 0 856 0 1 610
box 0 0 64 200
use AND2X2  _66_
timestamp 1656222261
transform -1 0 920 0 1 610
box 0 0 64 200
use XOR2X1  _65_
timestamp 1656222261
transform -1 0 1032 0 1 610
box 0 0 112 200
use AND2X2  _68_
timestamp 1656222261
transform -1 0 1096 0 1 610
box 0 0 64 200
use XOR2X1  _67_
timestamp 1656222261
transform -1 0 1208 0 1 610
box 0 0 112 200
use OR2X2  _33_
timestamp 1656222261
transform -1 0 1272 0 1 610
box 0 0 64 200
use AND2X2  _35_
timestamp 1656222261
transform -1 0 1336 0 1 610
box 0 0 64 200
use XOR2X1  _34_
timestamp 1656222261
transform -1 0 1448 0 1 610
box 0 0 112 200
use AND2X2  _37_
timestamp 1656222261
transform -1 0 1512 0 1 610
box 0 0 64 200
use XOR2X1  _36_
timestamp 1656222261
transform -1 0 1624 0 1 610
box 0 0 112 200
use OR2X2  _28_
timestamp 1656222261
transform -1 0 1688 0 1 610
box 0 0 64 200
use XOR2X1  _31_
timestamp 1656222261
transform 1 0 1688 0 1 610
box 0 0 112 200
use DFFSR  _12_
timestamp 1656222261
transform 1 0 1800 0 1 610
box 0 0 352 200
use FILL  FILL32280x9150
timestamp 1656222261
transform 1 0 2152 0 1 610
box 0 0 16 200
use AND2X2  _93_
timestamp 1656222261
transform 1 0 8 0 -1 610
box 0 0 64 200
use AND2X2  _135_
timestamp 1656222261
transform -1 0 136 0 -1 610
box 0 0 64 200
use XOR2X1  _144_
timestamp 1656222261
transform -1 0 248 0 -1 610
box 0 0 112 200
use AND2X2  _145_
timestamp 1656222261
transform 1 0 248 0 -1 610
box 0 0 64 200
use OR2X2  _143_
timestamp 1656222261
transform 1 0 312 0 -1 610
box 0 0 64 200
use AND2X2  _147_
timestamp 1656222261
transform -1 0 440 0 -1 610
box 0 0 64 200
use XOR2X1  _146_
timestamp 1656222261
transform -1 0 552 0 -1 610
box 0 0 112 200
use OR2X2  _109_
timestamp 1656222261
transform -1 0 616 0 -1 610
box 0 0 64 200
use XOR2X1  _39_
timestamp 1656222261
transform 1 0 616 0 -1 610
box 0 0 112 200
use AND2X2  _40_
timestamp 1656222261
transform 1 0 728 0 -1 610
box 0 0 64 200
use XOR2X1  _72_
timestamp 1656222261
transform -1 0 904 0 -1 610
box 0 0 112 200
use BUFX2  _4_
timestamp 1656222261
transform 1 0 904 0 -1 610
box 0 0 48 200
use OR2X2  _38_
timestamp 1656222261
transform 1 0 952 0 -1 610
box 0 0 64 200
use AND2X2  _42_
timestamp 1656222261
transform -1 0 1080 0 -1 610
box 0 0 64 200
use XOR2X1  _41_
timestamp 1656222261
transform -1 0 1192 0 -1 610
box 0 0 112 200
use DFFSR  _14_
timestamp 1656222261
transform -1 0 1544 0 -1 610
box 0 0 352 200
use BUFX2  BUFX2_insert1
timestamp 1656222261
transform -1 0 1592 0 -1 610
box 0 0 48 200
use BUFX2  BUFX2_insert3
timestamp 1656222261
transform -1 0 1640 0 -1 610
box 0 0 48 200
use AND2X2  _32_
timestamp 1656222261
transform -1 0 1704 0 -1 610
box 0 0 64 200
use DFFSR  _17_
timestamp 1656222261
transform -1 0 2056 0 -1 610
box 0 0 352 200
use XOR2X1  _29_
timestamp 1656222261
transform 1 0 2056 0 -1 610
box 0 0 112 200
use XOR2X1  _149_
timestamp 1656222261
transform -1 0 120 0 1 210
box 0 0 112 200
use AND2X2  _150_
timestamp 1656222261
transform 1 0 120 0 1 210
box 0 0 64 200
use AND2X2  _152_
timestamp 1656222261
transform -1 0 248 0 1 210
box 0 0 64 200
use XOR2X1  _151_
timestamp 1656222261
transform -1 0 360 0 1 210
box 0 0 112 200
use XOR2X1  _115_
timestamp 1656222261
transform -1 0 472 0 1 210
box 0 0 112 200
use AND2X2  _116_
timestamp 1656222261
transform 1 0 472 0 1 210
box 0 0 64 200
use AND2X2  _118_
timestamp 1656222261
transform -1 0 600 0 1 210
box 0 0 64 200
use XOR2X1  _117_
timestamp 1656222261
transform -1 0 712 0 1 210
box 0 0 112 200
use XOR2X1  _70_
timestamp 1656222261
transform 1 0 712 0 1 210
box 0 0 112 200
use AND2X2  _71_
timestamp 1656222261
transform 1 0 824 0 1 210
box 0 0 64 200
use AND2X2  _73_
timestamp 1656222261
transform 1 0 888 0 1 210
box 0 0 64 200
use OR2X2  _69_
timestamp 1656222261
transform 1 0 952 0 1 210
box 0 0 64 200
use XOR2X1  _46_
timestamp 1656222261
transform 1 0 1016 0 1 210
box 0 0 112 200
use AND2X2  _47_
timestamp 1656222261
transform 1 0 1128 0 1 210
box 0 0 64 200
use XOR2X1  _44_
timestamp 1656222261
transform -1 0 1304 0 1 210
box 0 0 112 200
use AND2X2  _45_
timestamp 1656222261
transform 1 0 1304 0 1 210
box 0 0 64 200
use OR2X2  _43_
timestamp 1656222261
transform 1 0 1368 0 1 210
box 0 0 64 200
use XOR2X1  _82_
timestamp 1656222261
transform 1 0 1432 0 1 210
box 0 0 112 200
use XOR2X1  _49_
timestamp 1656222261
transform 1 0 1544 0 1 210
box 0 0 112 200
use AND2X2  _50_
timestamp 1656222261
transform 1 0 1656 0 1 210
box 0 0 64 200
use XOR2X1  _51_
timestamp 1656222261
transform 1 0 1720 0 1 210
box 0 0 112 200
use AND2X2  _52_
timestamp 1656222261
transform 1 0 1832 0 1 210
box 0 0 64 200
use OR2X2  _48_
timestamp 1656222261
transform 1 0 1896 0 1 210
box 0 0 64 200
use XOR2X1  _53_
timestamp 1656222261
transform -1 0 2072 0 1 210
box 0 0 112 200
use BUFX2  _3_
timestamp 1656222261
transform 1 0 2072 0 1 210
box 0 0 48 200
use BUFX2  _7_
timestamp 1656222261
transform 1 0 2120 0 1 210
box 0 0 48 200
use XOR2X1  _120_
timestamp 1656222261
transform 1 0 8 0 -1 210
box 0 0 112 200
use OR2X2  _148_
timestamp 1656222261
transform -1 0 184 0 -1 210
box 0 0 64 200
use AND2X2  _121_
timestamp 1656222261
transform 1 0 184 0 -1 210
box 0 0 64 200
use OR2X2  _119_
timestamp 1656222261
transform 1 0 248 0 -1 210
box 0 0 64 200
use AND2X2  _123_
timestamp 1656222261
transform -1 0 376 0 -1 210
box 0 0 64 200
use XOR2X1  _122_
timestamp 1656222261
transform -1 0 488 0 -1 210
box 0 0 112 200
use OR2X2  _114_
timestamp 1656222261
transform -1 0 552 0 -1 210
box 0 0 64 200
use BUFX2  _5_
timestamp 1656222261
transform -1 0 600 0 -1 210
box 0 0 48 200
use XOR2X1  _75_
timestamp 1656222261
transform -1 0 712 0 -1 210
box 0 0 112 200
use BUFX2  _6_
timestamp 1656222261
transform -1 0 760 0 -1 210
box 0 0 48 200
use AND2X2  _76_
timestamp 1656222261
transform 1 0 760 0 -1 210
box 0 0 64 200
use DFFSR  _15_
timestamp 1656222261
transform -1 0 1176 0 -1 210
box 0 0 352 200
use XOR2X1  _77_
timestamp 1656222261
transform -1 0 1288 0 -1 210
box 0 0 112 200
use AND2X2  _78_
timestamp 1656222261
transform 1 0 1288 0 -1 210
box 0 0 64 200
use OR2X2  _74_
timestamp 1656222261
transform 1 0 1352 0 -1 210
box 0 0 64 200
use XOR2X1  _80_
timestamp 1656222261
transform -1 0 1528 0 -1 210
box 0 0 112 200
use AND2X2  _83_
timestamp 1656222261
transform 1 0 1528 0 -1 210
box 0 0 64 200
use AND2X2  _81_
timestamp 1656222261
transform 1 0 1592 0 -1 210
box 0 0 64 200
use OR2X2  _79_
timestamp 1656222261
transform 1 0 1656 0 -1 210
box 0 0 64 200
use AND2X2  _30_
timestamp 1656222261
transform -1 0 1784 0 -1 210
box 0 0 64 200
use DFFSR  _16_
timestamp 1656222261
transform 1 0 1784 0 -1 210
box 0 0 352 200
use FILL  FILL32040x150
timestamp 1656222261
transform -1 0 2152 0 -1 210
box 0 0 16 200
use FILL  FILL32280x150
timestamp 1656222261
transform -1 0 2168 0 -1 210
box 0 0 16 200
<< labels >>
flabel metal1 2178 4 2242 4 7 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 -66 4 -2 4 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal2 973 1457 979 1463 3 FreeSans 16 90 0 0 clk
port 2 nsew
flabel metal3 2203 895 2213 905 3 FreeSans 16 0 0 0 f[8]
port 3 nsew
flabel metal3 2203 295 2213 305 3 FreeSans 16 0 0 0 f[7]
port 4 nsew
flabel metal2 733 -23 739 -17 7 FreeSans 16 270 0 0 f[6]
port 5 nsew
flabel metal2 573 -23 579 -17 7 FreeSans 16 270 0 0 f[5]
port 6 nsew
flabel metal2 925 -23 931 -17 7 FreeSans 16 270 0 0 f[4]
port 7 nsew
flabel metal3 2203 335 2213 345 3 FreeSans 16 0 0 0 f[3]
port 8 nsew
flabel metal3 2203 1295 2213 1305 3 FreeSans 16 0 0 0 f[2]
port 9 nsew
flabel metal2 1341 1457 1347 1463 3 FreeSans 16 90 0 0 f[1]
port 10 nsew
flabel metal2 765 1457 771 1463 3 FreeSans 16 90 0 0 f[0]
port 11 nsew
flabel metal3 -37 715 -27 725 7 FreeSans 16 0 0 0 i[3]
port 12 nsew
flabel metal3 -37 515 -27 525 7 FreeSans 16 0 0 0 i[2]
port 13 nsew
flabel metal3 -37 915 -27 925 7 FreeSans 16 0 0 0 i[1]
port 14 nsew
flabel metal2 509 1457 515 1463 3 FreeSans 16 90 0 0 i[0]
port 15 nsew
flabel metal3 -37 555 -27 565 7 FreeSans 16 0 0 0 j[3]
port 16 nsew
flabel metal3 -37 1295 -27 1305 7 FreeSans 16 0 0 0 j[2]
port 17 nsew
flabel metal2 541 1457 547 1463 3 FreeSans 16 90 0 0 j[1]
port 18 nsew
flabel metal2 461 1457 467 1463 3 FreeSans 16 90 0 0 j[0]
port 19 nsew
flabel metal2 1069 1457 1075 1463 3 FreeSans 16 90 0 0 rst
port 20 nsew
<< end >>
